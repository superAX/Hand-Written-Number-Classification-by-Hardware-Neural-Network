`timescale 1 ns/10 ps
module Image_Classifier ( 
  input clk, 
  input GlobalReset, 
  input Input_Valid,
  input [18:0] Wgt_0_0, // sfix19_En18 
  input [18:0] Wgt_0_1, // sfix19_En18 
  input [18:0] Wgt_0_2, // sfix19_En18 
  input [18:0] Wgt_0_3, // sfix19_En18 
  input [18:0] Wgt_0_4, // sfix19_En18 
  input [18:0] Wgt_0_5, // sfix19_En18 
  input [18:0] Wgt_0_6, // sfix19_En18 
  input [18:0] Wgt_0_7, // sfix19_En18 
  input [18:0] Wgt_0_8, // sfix19_En18 
  input [18:0] Wgt_0_9, // sfix19_En18 
  input [18:0] Wgt_0_10, // sfix19_En18 
  input [18:0] Wgt_0_11, // sfix19_En18 
  input [18:0] Wgt_0_12, // sfix19_En18 
  input [18:0] Wgt_0_13, // sfix19_En18 
  input [18:0] Wgt_0_14, // sfix19_En18 
  input [18:0] Wgt_0_15, // sfix19_En18 
  input [18:0] Wgt_0_16, // sfix19_En18 
  input [18:0] Wgt_0_17, // sfix19_En18 
  input [18:0] Wgt_0_18, // sfix19_En18 
  input [18:0] Wgt_0_19, // sfix19_En18 
  input [18:0] Wgt_0_20, // sfix19_En18 
  input [18:0] Wgt_0_21, // sfix19_En18 
  input [18:0] Wgt_0_22, // sfix19_En18 
  input [18:0] Wgt_0_23, // sfix19_En18 
  input [18:0] Wgt_0_24, // sfix19_En18 
  input [18:0] Wgt_0_25, // sfix19_En18 
  input [18:0] Wgt_0_26, // sfix19_En18 
  input [18:0] Wgt_0_27, // sfix19_En18 
  input [18:0] Wgt_0_28, // sfix19_En18 
  input [18:0] Wgt_0_29, // sfix19_En18 
  input [18:0] Wgt_0_30, // sfix19_En18 
  input [18:0] Wgt_0_31, // sfix19_En18 
  input [18:0] Wgt_0_32, // sfix19_En18 
  input [18:0] Wgt_0_33, // sfix19_En18 
  input [18:0] Wgt_0_34, // sfix19_En18 
  input [18:0] Wgt_0_35, // sfix19_En18 
  input [18:0] Wgt_0_36, // sfix19_En18 
  input [18:0] Wgt_0_37, // sfix19_En18 
  input [18:0] Wgt_0_38, // sfix19_En18 
  input [18:0] Wgt_0_39, // sfix19_En18 
  input [18:0] Wgt_0_40, // sfix19_En18 
  input [18:0] Wgt_0_41, // sfix19_En18 
  input [18:0] Wgt_0_42, // sfix19_En18 
  input [18:0] Wgt_0_43, // sfix19_En18 
  input [18:0] Wgt_0_44, // sfix19_En18 
  input [18:0] Wgt_0_45, // sfix19_En18 
  input [18:0] Wgt_0_46, // sfix19_En18 
  input [18:0] Wgt_0_47, // sfix19_En18 
  input [18:0] Wgt_0_48, // sfix19_En18 
  input [18:0] Wgt_0_49, // sfix19_En18 
  input [18:0] Wgt_0_50, // sfix19_En18 
  input [18:0] Wgt_0_51, // sfix19_En18 
  input [18:0] Wgt_0_52, // sfix19_En18 
  input [18:0] Wgt_0_53, // sfix19_En18 
  input [18:0] Wgt_0_54, // sfix19_En18 
  input [18:0] Wgt_0_55, // sfix19_En18 
  input [18:0] Wgt_0_56, // sfix19_En18 
  input [18:0] Wgt_0_57, // sfix19_En18 
  input [18:0] Wgt_0_58, // sfix19_En18 
  input [18:0] Wgt_0_59, // sfix19_En18 
  input [18:0] Wgt_0_60, // sfix19_En18 
  input [18:0] Wgt_0_61, // sfix19_En18 
  input [18:0] Wgt_0_62, // sfix19_En18 
  input [18:0] Wgt_0_63, // sfix19_En18 
  input [18:0] Wgt_0_64, // sfix19_En18 
  input [18:0] Wgt_0_65, // sfix19_En18 
  input [18:0] Wgt_0_66, // sfix19_En18 
  input [18:0] Wgt_0_67, // sfix19_En18 
  input [18:0] Wgt_0_68, // sfix19_En18 
  input [18:0] Wgt_0_69, // sfix19_En18 
  input [18:0] Wgt_0_70, // sfix19_En18 
  input [18:0] Wgt_0_71, // sfix19_En18 
  input [18:0] Wgt_0_72, // sfix19_En18 
  input [18:0] Wgt_0_73, // sfix19_En18 
  input [18:0] Wgt_0_74, // sfix19_En18 
  input [18:0] Wgt_0_75, // sfix19_En18 
  input [18:0] Wgt_0_76, // sfix19_En18 
  input [18:0] Wgt_0_77, // sfix19_En18 
  input [18:0] Wgt_0_78, // sfix19_En18 
  input [18:0] Wgt_0_79, // sfix19_En18 
  input [18:0] Wgt_0_80, // sfix19_En18 
  input [18:0] Wgt_0_81, // sfix19_En18 
  input [18:0] Wgt_0_82, // sfix19_En18 
  input [18:0] Wgt_0_83, // sfix19_En18 
  input [18:0] Wgt_0_84, // sfix19_En18 
  input [18:0] Wgt_0_85, // sfix19_En18 
  input [18:0] Wgt_0_86, // sfix19_En18 
  input [18:0] Wgt_0_87, // sfix19_En18 
  input [18:0] Wgt_0_88, // sfix19_En18 
  input [18:0] Wgt_0_89, // sfix19_En18 
  input [18:0] Wgt_0_90, // sfix19_En18 
  input [18:0] Wgt_0_91, // sfix19_En18 
  input [18:0] Wgt_0_92, // sfix19_En18 
  input [18:0] Wgt_0_93, // sfix19_En18 
  input [18:0] Wgt_0_94, // sfix19_En18 
  input [18:0] Wgt_0_95, // sfix19_En18 
  input [18:0] Wgt_0_96, // sfix19_En18 
  input [18:0] Wgt_0_97, // sfix19_En18 
  input [18:0] Wgt_0_98, // sfix19_En18 
  input [18:0] Wgt_0_99, // sfix19_En18 
  input [18:0] Wgt_0_100, // sfix19_En18 
  input [18:0] Wgt_0_101, // sfix19_En18 
  input [18:0] Wgt_0_102, // sfix19_En18 
  input [18:0] Wgt_0_103, // sfix19_En18 
  input [18:0] Wgt_0_104, // sfix19_En18 
  input [18:0] Wgt_0_105, // sfix19_En18 
  input [18:0] Wgt_0_106, // sfix19_En18 
  input [18:0] Wgt_0_107, // sfix19_En18 
  input [18:0] Wgt_0_108, // sfix19_En18 
  input [18:0] Wgt_0_109, // sfix19_En18 
  input [18:0] Wgt_0_110, // sfix19_En18 
  input [18:0] Wgt_0_111, // sfix19_En18 
  input [18:0] Wgt_0_112, // sfix19_En18 
  input [18:0] Wgt_0_113, // sfix19_En18 
  input [18:0] Wgt_0_114, // sfix19_En18 
  input [18:0] Wgt_0_115, // sfix19_En18 
  input [18:0] Wgt_0_116, // sfix19_En18 
  input [18:0] Wgt_0_117, // sfix19_En18 
  input [18:0] Wgt_0_118, // sfix19_En18 
  input [18:0] Wgt_0_119, // sfix19_En18 
  input [18:0] Wgt_0_120, // sfix19_En18 
  input [18:0] Wgt_0_121, // sfix19_En18 
  input [18:0] Wgt_0_122, // sfix19_En18 
  input [18:0] Wgt_0_123, // sfix19_En18 
  input [18:0] Wgt_0_124, // sfix19_En18 
  input [18:0] Wgt_0_125, // sfix19_En18 
  input [18:0] Wgt_0_126, // sfix19_En18 
  input [18:0] Wgt_0_127, // sfix19_En18 
  input [18:0] Wgt_0_128, // sfix19_En18 
  input [18:0] Wgt_0_129, // sfix19_En18 
  input [18:0] Wgt_0_130, // sfix19_En18 
  input [18:0] Wgt_0_131, // sfix19_En18 
  input [18:0] Wgt_0_132, // sfix19_En18 
  input [18:0] Wgt_0_133, // sfix19_En18 
  input [18:0] Wgt_0_134, // sfix19_En18 
  input [18:0] Wgt_0_135, // sfix19_En18 
  input [18:0] Wgt_0_136, // sfix19_En18 
  input [18:0] Wgt_0_137, // sfix19_En18 
  input [18:0] Wgt_0_138, // sfix19_En18 
  input [18:0] Wgt_0_139, // sfix19_En18 
  input [18:0] Wgt_0_140, // sfix19_En18 
  input [18:0] Wgt_0_141, // sfix19_En18 
  input [18:0] Wgt_0_142, // sfix19_En18 
  input [18:0] Wgt_0_143, // sfix19_En18 
  input [18:0] Wgt_0_144, // sfix19_En18 
  input [18:0] Wgt_0_145, // sfix19_En18 
  input [18:0] Wgt_0_146, // sfix19_En18 
  input [18:0] Wgt_0_147, // sfix19_En18 
  input [18:0] Wgt_0_148, // sfix19_En18 
  input [18:0] Wgt_0_149, // sfix19_En18 
  input [18:0] Wgt_0_150, // sfix19_En18 
  input [18:0] Wgt_0_151, // sfix19_En18 
  input [18:0] Wgt_0_152, // sfix19_En18 
  input [18:0] Wgt_0_153, // sfix19_En18 
  input [18:0] Wgt_0_154, // sfix19_En18 
  input [18:0] Wgt_0_155, // sfix19_En18 
  input [18:0] Wgt_0_156, // sfix19_En18 
  input [18:0] Wgt_0_157, // sfix19_En18 
  input [18:0] Wgt_0_158, // sfix19_En18 
  input [18:0] Wgt_0_159, // sfix19_En18 
  input [18:0] Wgt_0_160, // sfix19_En18 
  input [18:0] Wgt_0_161, // sfix19_En18 
  input [18:0] Wgt_0_162, // sfix19_En18 
  input [18:0] Wgt_0_163, // sfix19_En18 
  input [18:0] Wgt_0_164, // sfix19_En18 
  input [18:0] Wgt_0_165, // sfix19_En18 
  input [18:0] Wgt_0_166, // sfix19_En18 
  input [18:0] Wgt_0_167, // sfix19_En18 
  input [18:0] Wgt_0_168, // sfix19_En18 
  input [18:0] Wgt_0_169, // sfix19_En18 
  input [18:0] Wgt_0_170, // sfix19_En18 
  input [18:0] Wgt_0_171, // sfix19_En18 
  input [18:0] Wgt_0_172, // sfix19_En18 
  input [18:0] Wgt_0_173, // sfix19_En18 
  input [18:0] Wgt_0_174, // sfix19_En18 
  input [18:0] Wgt_0_175, // sfix19_En18 
  input [18:0] Wgt_0_176, // sfix19_En18 
  input [18:0] Wgt_0_177, // sfix19_En18 
  input [18:0] Wgt_0_178, // sfix19_En18 
  input [18:0] Wgt_0_179, // sfix19_En18 
  input [18:0] Wgt_0_180, // sfix19_En18 
  input [18:0] Wgt_0_181, // sfix19_En18 
  input [18:0] Wgt_0_182, // sfix19_En18 
  input [18:0] Wgt_0_183, // sfix19_En18 
  input [18:0] Wgt_0_184, // sfix19_En18 
  input [18:0] Wgt_0_185, // sfix19_En18 
  input [18:0] Wgt_0_186, // sfix19_En18 
  input [18:0] Wgt_0_187, // sfix19_En18 
  input [18:0] Wgt_0_188, // sfix19_En18 
  input [18:0] Wgt_0_189, // sfix19_En18 
  input [18:0] Wgt_0_190, // sfix19_En18 
  input [18:0] Wgt_0_191, // sfix19_En18 
  input [18:0] Wgt_0_192, // sfix19_En18 
  input [18:0] Wgt_0_193, // sfix19_En18 
  input [18:0] Wgt_0_194, // sfix19_En18 
  input [18:0] Wgt_0_195, // sfix19_En18 
  input [18:0] Wgt_0_196, // sfix19_En18 
  input [18:0] Wgt_0_197, // sfix19_En18 
  input [18:0] Wgt_0_198, // sfix19_En18 
  input [18:0] Wgt_0_199, // sfix19_En18 
  input [18:0] Wgt_0_200, // sfix19_En18 
  input [18:0] Wgt_0_201, // sfix19_En18 
  input [18:0] Wgt_0_202, // sfix19_En18 
  input [18:0] Wgt_0_203, // sfix19_En18 
  input [18:0] Wgt_0_204, // sfix19_En18 
  input [18:0] Wgt_0_205, // sfix19_En18 
  input [18:0] Wgt_0_206, // sfix19_En18 
  input [18:0] Wgt_0_207, // sfix19_En18 
  input [18:0] Wgt_0_208, // sfix19_En18 
  input [18:0] Wgt_0_209, // sfix19_En18 
  input [18:0] Wgt_0_210, // sfix19_En18 
  input [18:0] Wgt_0_211, // sfix19_En18 
  input [18:0] Wgt_0_212, // sfix19_En18 
  input [18:0] Wgt_0_213, // sfix19_En18 
  input [18:0] Wgt_0_214, // sfix19_En18 
  input [18:0] Wgt_0_215, // sfix19_En18 
  input [18:0] Wgt_0_216, // sfix19_En18 
  input [18:0] Wgt_0_217, // sfix19_En18 
  input [18:0] Wgt_0_218, // sfix19_En18 
  input [18:0] Wgt_0_219, // sfix19_En18 
  input [18:0] Wgt_0_220, // sfix19_En18 
  input [18:0] Wgt_0_221, // sfix19_En18 
  input [18:0] Wgt_0_222, // sfix19_En18 
  input [18:0] Wgt_0_223, // sfix19_En18 
  input [18:0] Wgt_0_224, // sfix19_En18 
  input [18:0] Wgt_0_225, // sfix19_En18 
  input [18:0] Wgt_0_226, // sfix19_En18 
  input [18:0] Wgt_0_227, // sfix19_En18 
  input [18:0] Wgt_0_228, // sfix19_En18 
  input [18:0] Wgt_0_229, // sfix19_En18 
  input [18:0] Wgt_0_230, // sfix19_En18 
  input [18:0] Wgt_0_231, // sfix19_En18 
  input [18:0] Wgt_0_232, // sfix19_En18 
  input [18:0] Wgt_0_233, // sfix19_En18 
  input [18:0] Wgt_0_234, // sfix19_En18 
  input [18:0] Wgt_0_235, // sfix19_En18 
  input [18:0] Wgt_0_236, // sfix19_En18 
  input [18:0] Wgt_0_237, // sfix19_En18 
  input [18:0] Wgt_0_238, // sfix19_En18 
  input [18:0] Wgt_0_239, // sfix19_En18 
  input [18:0] Wgt_0_240, // sfix19_En18 
  input [18:0] Wgt_0_241, // sfix19_En18 
  input [18:0] Wgt_0_242, // sfix19_En18 
  input [18:0] Wgt_0_243, // sfix19_En18 
  input [18:0] Wgt_0_244, // sfix19_En18 
  input [18:0] Wgt_0_245, // sfix19_En18 
  input [18:0] Wgt_0_246, // sfix19_En18 
  input [18:0] Wgt_0_247, // sfix19_En18 
  input [18:0] Wgt_0_248, // sfix19_En18 
  input [18:0] Wgt_0_249, // sfix19_En18 
  input [18:0] Wgt_0_250, // sfix19_En18 
  input [18:0] Wgt_0_251, // sfix19_En18 
  input [18:0] Wgt_0_252, // sfix19_En18 
  input [18:0] Wgt_0_253, // sfix19_En18 
  input [18:0] Wgt_0_254, // sfix19_En18 
  input [18:0] Wgt_0_255, // sfix19_En18 
  input [18:0] Wgt_0_256, // sfix19_En18 
  input [18:0] Wgt_0_257, // sfix19_En18 
  input [18:0] Wgt_0_258, // sfix19_En18 
  input [18:0] Wgt_0_259, // sfix19_En18 
  input [18:0] Wgt_0_260, // sfix19_En18 
  input [18:0] Wgt_0_261, // sfix19_En18 
  input [18:0] Wgt_0_262, // sfix19_En18 
  input [18:0] Wgt_0_263, // sfix19_En18 
  input [18:0] Wgt_0_264, // sfix19_En18 
  input [18:0] Wgt_0_265, // sfix19_En18 
  input [18:0] Wgt_0_266, // sfix19_En18 
  input [18:0] Wgt_0_267, // sfix19_En18 
  input [18:0] Wgt_0_268, // sfix19_En18 
  input [18:0] Wgt_0_269, // sfix19_En18 
  input [18:0] Wgt_0_270, // sfix19_En18 
  input [18:0] Wgt_0_271, // sfix19_En18 
  input [18:0] Wgt_0_272, // sfix19_En18 
  input [18:0] Wgt_0_273, // sfix19_En18 
  input [18:0] Wgt_0_274, // sfix19_En18 
  input [18:0] Wgt_0_275, // sfix19_En18 
  input [18:0] Wgt_0_276, // sfix19_En18 
  input [18:0] Wgt_0_277, // sfix19_En18 
  input [18:0] Wgt_0_278, // sfix19_En18 
  input [18:0] Wgt_0_279, // sfix19_En18 
  input [18:0] Wgt_0_280, // sfix19_En18 
  input [18:0] Wgt_0_281, // sfix19_En18 
  input [18:0] Wgt_0_282, // sfix19_En18 
  input [18:0] Wgt_0_283, // sfix19_En18 
  input [18:0] Wgt_0_284, // sfix19_En18 
  input [18:0] Wgt_0_285, // sfix19_En18 
  input [18:0] Wgt_0_286, // sfix19_En18 
  input [18:0] Wgt_0_287, // sfix19_En18 
  input [18:0] Wgt_0_288, // sfix19_En18 
  input [18:0] Wgt_0_289, // sfix19_En18 
  input [18:0] Wgt_0_290, // sfix19_En18 
  input [18:0] Wgt_0_291, // sfix19_En18 
  input [18:0] Wgt_0_292, // sfix19_En18 
  input [18:0] Wgt_0_293, // sfix19_En18 
  input [18:0] Wgt_0_294, // sfix19_En18 
  input [18:0] Wgt_0_295, // sfix19_En18 
  input [18:0] Wgt_0_296, // sfix19_En18 
  input [18:0] Wgt_0_297, // sfix19_En18 
  input [18:0] Wgt_0_298, // sfix19_En18 
  input [18:0] Wgt_0_299, // sfix19_En18 
  input [18:0] Wgt_0_300, // sfix19_En18 
  input [18:0] Wgt_0_301, // sfix19_En18 
  input [18:0] Wgt_0_302, // sfix19_En18 
  input [18:0] Wgt_0_303, // sfix19_En18 
  input [18:0] Wgt_0_304, // sfix19_En18 
  input [18:0] Wgt_0_305, // sfix19_En18 
  input [18:0] Wgt_0_306, // sfix19_En18 
  input [18:0] Wgt_0_307, // sfix19_En18 
  input [18:0] Wgt_0_308, // sfix19_En18 
  input [18:0] Wgt_0_309, // sfix19_En18 
  input [18:0] Wgt_0_310, // sfix19_En18 
  input [18:0] Wgt_0_311, // sfix19_En18 
  input [18:0] Wgt_0_312, // sfix19_En18 
  input [18:0] Wgt_0_313, // sfix19_En18 
  input [18:0] Wgt_0_314, // sfix19_En18 
  input [18:0] Wgt_0_315, // sfix19_En18 
  input [18:0] Wgt_0_316, // sfix19_En18 
  input [18:0] Wgt_0_317, // sfix19_En18 
  input [18:0] Wgt_0_318, // sfix19_En18 
  input [18:0] Wgt_0_319, // sfix19_En18 
  input [18:0] Wgt_0_320, // sfix19_En18 
  input [18:0] Wgt_0_321, // sfix19_En18 
  input [18:0] Wgt_0_322, // sfix19_En18 
  input [18:0] Wgt_0_323, // sfix19_En18 
  input [18:0] Wgt_0_324, // sfix19_En18 
  input [18:0] Wgt_0_325, // sfix19_En18 
  input [18:0] Wgt_0_326, // sfix19_En18 
  input [18:0] Wgt_0_327, // sfix19_En18 
  input [18:0] Wgt_0_328, // sfix19_En18 
  input [18:0] Wgt_0_329, // sfix19_En18 
  input [18:0] Wgt_0_330, // sfix19_En18 
  input [18:0] Wgt_0_331, // sfix19_En18 
  input [18:0] Wgt_0_332, // sfix19_En18 
  input [18:0] Wgt_0_333, // sfix19_En18 
  input [18:0] Wgt_0_334, // sfix19_En18 
  input [18:0] Wgt_0_335, // sfix19_En18 
  input [18:0] Wgt_0_336, // sfix19_En18 
  input [18:0] Wgt_0_337, // sfix19_En18 
  input [18:0] Wgt_0_338, // sfix19_En18 
  input [18:0] Wgt_0_339, // sfix19_En18 
  input [18:0] Wgt_0_340, // sfix19_En18 
  input [18:0] Wgt_0_341, // sfix19_En18 
  input [18:0] Wgt_0_342, // sfix19_En18 
  input [18:0] Wgt_0_343, // sfix19_En18 
  input [18:0] Wgt_0_344, // sfix19_En18 
  input [18:0] Wgt_0_345, // sfix19_En18 
  input [18:0] Wgt_0_346, // sfix19_En18 
  input [18:0] Wgt_0_347, // sfix19_En18 
  input [18:0] Wgt_0_348, // sfix19_En18 
  input [18:0] Wgt_0_349, // sfix19_En18 
  input [18:0] Wgt_0_350, // sfix19_En18 
  input [18:0] Wgt_0_351, // sfix19_En18 
  input [18:0] Wgt_0_352, // sfix19_En18 
  input [18:0] Wgt_0_353, // sfix19_En18 
  input [18:0] Wgt_0_354, // sfix19_En18 
  input [18:0] Wgt_0_355, // sfix19_En18 
  input [18:0] Wgt_0_356, // sfix19_En18 
  input [18:0] Wgt_0_357, // sfix19_En18 
  input [18:0] Wgt_0_358, // sfix19_En18 
  input [18:0] Wgt_0_359, // sfix19_En18 
  input [18:0] Wgt_0_360, // sfix19_En18 
  input [18:0] Wgt_0_361, // sfix19_En18 
  input [18:0] Wgt_0_362, // sfix19_En18 
  input [18:0] Wgt_0_363, // sfix19_En18 
  input [18:0] Wgt_0_364, // sfix19_En18 
  input [18:0] Wgt_0_365, // sfix19_En18 
  input [18:0] Wgt_0_366, // sfix19_En18 
  input [18:0] Wgt_0_367, // sfix19_En18 
  input [18:0] Wgt_0_368, // sfix19_En18 
  input [18:0] Wgt_0_369, // sfix19_En18 
  input [18:0] Wgt_0_370, // sfix19_En18 
  input [18:0] Wgt_0_371, // sfix19_En18 
  input [18:0] Wgt_0_372, // sfix19_En18 
  input [18:0] Wgt_0_373, // sfix19_En18 
  input [18:0] Wgt_0_374, // sfix19_En18 
  input [18:0] Wgt_0_375, // sfix19_En18 
  input [18:0] Wgt_0_376, // sfix19_En18 
  input [18:0] Wgt_0_377, // sfix19_En18 
  input [18:0] Wgt_0_378, // sfix19_En18 
  input [18:0] Wgt_0_379, // sfix19_En18 
  input [18:0] Wgt_0_380, // sfix19_En18 
  input [18:0] Wgt_0_381, // sfix19_En18 
  input [18:0] Wgt_0_382, // sfix19_En18 
  input [18:0] Wgt_0_383, // sfix19_En18 
  input [18:0] Wgt_0_384, // sfix19_En18 
  input [18:0] Wgt_0_385, // sfix19_En18 
  input [18:0] Wgt_0_386, // sfix19_En18 
  input [18:0] Wgt_0_387, // sfix19_En18 
  input [18:0] Wgt_0_388, // sfix19_En18 
  input [18:0] Wgt_0_389, // sfix19_En18 
  input [18:0] Wgt_0_390, // sfix19_En18 
  input [18:0] Wgt_0_391, // sfix19_En18 
  input [18:0] Wgt_0_392, // sfix19_En18 
  input [18:0] Wgt_0_393, // sfix19_En18 
  input [18:0] Wgt_0_394, // sfix19_En18 
  input [18:0] Wgt_0_395, // sfix19_En18 
  input [18:0] Wgt_0_396, // sfix19_En18 
  input [18:0] Wgt_0_397, // sfix19_En18 
  input [18:0] Wgt_0_398, // sfix19_En18 
  input [18:0] Wgt_0_399, // sfix19_En18 
  input [18:0] Wgt_0_400, // sfix19_En18 
  input [18:0] Wgt_0_401, // sfix19_En18 
  input [18:0] Wgt_0_402, // sfix19_En18 
  input [18:0] Wgt_0_403, // sfix19_En18 
  input [18:0] Wgt_0_404, // sfix19_En18 
  input [18:0] Wgt_0_405, // sfix19_En18 
  input [18:0] Wgt_0_406, // sfix19_En18 
  input [18:0] Wgt_0_407, // sfix19_En18 
  input [18:0] Wgt_0_408, // sfix19_En18 
  input [18:0] Wgt_0_409, // sfix19_En18 
  input [18:0] Wgt_0_410, // sfix19_En18 
  input [18:0] Wgt_0_411, // sfix19_En18 
  input [18:0] Wgt_0_412, // sfix19_En18 
  input [18:0] Wgt_0_413, // sfix19_En18 
  input [18:0] Wgt_0_414, // sfix19_En18 
  input [18:0] Wgt_0_415, // sfix19_En18 
  input [18:0] Wgt_0_416, // sfix19_En18 
  input [18:0] Wgt_0_417, // sfix19_En18 
  input [18:0] Wgt_0_418, // sfix19_En18 
  input [18:0] Wgt_0_419, // sfix19_En18 
  input [18:0] Wgt_0_420, // sfix19_En18 
  input [18:0] Wgt_0_421, // sfix19_En18 
  input [18:0] Wgt_0_422, // sfix19_En18 
  input [18:0] Wgt_0_423, // sfix19_En18 
  input [18:0] Wgt_0_424, // sfix19_En18 
  input [18:0] Wgt_0_425, // sfix19_En18 
  input [18:0] Wgt_0_426, // sfix19_En18 
  input [18:0] Wgt_0_427, // sfix19_En18 
  input [18:0] Wgt_0_428, // sfix19_En18 
  input [18:0] Wgt_0_429, // sfix19_En18 
  input [18:0] Wgt_0_430, // sfix19_En18 
  input [18:0] Wgt_0_431, // sfix19_En18 
  input [18:0] Wgt_0_432, // sfix19_En18 
  input [18:0] Wgt_0_433, // sfix19_En18 
  input [18:0] Wgt_0_434, // sfix19_En18 
  input [18:0] Wgt_0_435, // sfix19_En18 
  input [18:0] Wgt_0_436, // sfix19_En18 
  input [18:0] Wgt_0_437, // sfix19_En18 
  input [18:0] Wgt_0_438, // sfix19_En18 
  input [18:0] Wgt_0_439, // sfix19_En18 
  input [18:0] Wgt_0_440, // sfix19_En18 
  input [18:0] Wgt_0_441, // sfix19_En18 
  input [18:0] Wgt_0_442, // sfix19_En18 
  input [18:0] Wgt_0_443, // sfix19_En18 
  input [18:0] Wgt_0_444, // sfix19_En18 
  input [18:0] Wgt_0_445, // sfix19_En18 
  input [18:0] Wgt_0_446, // sfix19_En18 
  input [18:0] Wgt_0_447, // sfix19_En18 
  input [18:0] Wgt_0_448, // sfix19_En18 
  input [18:0] Wgt_0_449, // sfix19_En18 
  input [18:0] Wgt_0_450, // sfix19_En18 
  input [18:0] Wgt_0_451, // sfix19_En18 
  input [18:0] Wgt_0_452, // sfix19_En18 
  input [18:0] Wgt_0_453, // sfix19_En18 
  input [18:0] Wgt_0_454, // sfix19_En18 
  input [18:0] Wgt_0_455, // sfix19_En18 
  input [18:0] Wgt_0_456, // sfix19_En18 
  input [18:0] Wgt_0_457, // sfix19_En18 
  input [18:0] Wgt_0_458, // sfix19_En18 
  input [18:0] Wgt_0_459, // sfix19_En18 
  input [18:0] Wgt_0_460, // sfix19_En18 
  input [18:0] Wgt_0_461, // sfix19_En18 
  input [18:0] Wgt_0_462, // sfix19_En18 
  input [18:0] Wgt_0_463, // sfix19_En18 
  input [18:0] Wgt_0_464, // sfix19_En18 
  input [18:0] Wgt_0_465, // sfix19_En18 
  input [18:0] Wgt_0_466, // sfix19_En18 
  input [18:0] Wgt_0_467, // sfix19_En18 
  input [18:0] Wgt_0_468, // sfix19_En18 
  input [18:0] Wgt_0_469, // sfix19_En18 
  input [18:0] Wgt_0_470, // sfix19_En18 
  input [18:0] Wgt_0_471, // sfix19_En18 
  input [18:0] Wgt_0_472, // sfix19_En18 
  input [18:0] Wgt_0_473, // sfix19_En18 
  input [18:0] Wgt_0_474, // sfix19_En18 
  input [18:0] Wgt_0_475, // sfix19_En18 
  input [18:0] Wgt_0_476, // sfix19_En18 
  input [18:0] Wgt_0_477, // sfix19_En18 
  input [18:0] Wgt_0_478, // sfix19_En18 
  input [18:0] Wgt_0_479, // sfix19_En18 
  input [18:0] Wgt_0_480, // sfix19_En18 
  input [18:0] Wgt_0_481, // sfix19_En18 
  input [18:0] Wgt_0_482, // sfix19_En18 
  input [18:0] Wgt_0_483, // sfix19_En18 
  input [18:0] Wgt_0_484, // sfix19_En18 
  input [18:0] Wgt_0_485, // sfix19_En18 
  input [18:0] Wgt_0_486, // sfix19_En18 
  input [18:0] Wgt_0_487, // sfix19_En18 
  input [18:0] Wgt_0_488, // sfix19_En18 
  input [18:0] Wgt_0_489, // sfix19_En18 
  input [18:0] Wgt_0_490, // sfix19_En18 
  input [18:0] Wgt_0_491, // sfix19_En18 
  input [18:0] Wgt_0_492, // sfix19_En18 
  input [18:0] Wgt_0_493, // sfix19_En18 
  input [18:0] Wgt_0_494, // sfix19_En18 
  input [18:0] Wgt_0_495, // sfix19_En18 
  input [18:0] Wgt_0_496, // sfix19_En18 
  input [18:0] Wgt_0_497, // sfix19_En18 
  input [18:0] Wgt_0_498, // sfix19_En18 
  input [18:0] Wgt_0_499, // sfix19_En18 
  input [18:0] Wgt_0_500, // sfix19_En18 
  input [18:0] Wgt_0_501, // sfix19_En18 
  input [18:0] Wgt_0_502, // sfix19_En18 
  input [18:0] Wgt_0_503, // sfix19_En18 
  input [18:0] Wgt_0_504, // sfix19_En18 
  input [18:0] Wgt_0_505, // sfix19_En18 
  input [18:0] Wgt_0_506, // sfix19_En18 
  input [18:0] Wgt_0_507, // sfix19_En18 
  input [18:0] Wgt_0_508, // sfix19_En18 
  input [18:0] Wgt_0_509, // sfix19_En18 
  input [18:0] Wgt_0_510, // sfix19_En18 
  input [18:0] Wgt_0_511, // sfix19_En18 
  input [18:0] Wgt_0_512, // sfix19_En18 
  input [18:0] Wgt_0_513, // sfix19_En18 
  input [18:0] Wgt_0_514, // sfix19_En18 
  input [18:0] Wgt_0_515, // sfix19_En18 
  input [18:0] Wgt_0_516, // sfix19_En18 
  input [18:0] Wgt_0_517, // sfix19_En18 
  input [18:0] Wgt_0_518, // sfix19_En18 
  input [18:0] Wgt_0_519, // sfix19_En18 
  input [18:0] Wgt_0_520, // sfix19_En18 
  input [18:0] Wgt_0_521, // sfix19_En18 
  input [18:0] Wgt_0_522, // sfix19_En18 
  input [18:0] Wgt_0_523, // sfix19_En18 
  input [18:0] Wgt_0_524, // sfix19_En18 
  input [18:0] Wgt_0_525, // sfix19_En18 
  input [18:0] Wgt_0_526, // sfix19_En18 
  input [18:0] Wgt_0_527, // sfix19_En18 
  input [18:0] Wgt_0_528, // sfix19_En18 
  input [18:0] Wgt_0_529, // sfix19_En18 
  input [18:0] Wgt_0_530, // sfix19_En18 
  input [18:0] Wgt_0_531, // sfix19_En18 
  input [18:0] Wgt_0_532, // sfix19_En18 
  input [18:0] Wgt_0_533, // sfix19_En18 
  input [18:0] Wgt_0_534, // sfix19_En18 
  input [18:0] Wgt_0_535, // sfix19_En18 
  input [18:0] Wgt_0_536, // sfix19_En18 
  input [18:0] Wgt_0_537, // sfix19_En18 
  input [18:0] Wgt_0_538, // sfix19_En18 
  input [18:0] Wgt_0_539, // sfix19_En18 
  input [18:0] Wgt_0_540, // sfix19_En18 
  input [18:0] Wgt_0_541, // sfix19_En18 
  input [18:0] Wgt_0_542, // sfix19_En18 
  input [18:0] Wgt_0_543, // sfix19_En18 
  input [18:0] Wgt_0_544, // sfix19_En18 
  input [18:0] Wgt_0_545, // sfix19_En18 
  input [18:0] Wgt_0_546, // sfix19_En18 
  input [18:0] Wgt_0_547, // sfix19_En18 
  input [18:0] Wgt_0_548, // sfix19_En18 
  input [18:0] Wgt_0_549, // sfix19_En18 
  input [18:0] Wgt_0_550, // sfix19_En18 
  input [18:0] Wgt_0_551, // sfix19_En18 
  input [18:0] Wgt_0_552, // sfix19_En18 
  input [18:0] Wgt_0_553, // sfix19_En18 
  input [18:0] Wgt_0_554, // sfix19_En18 
  input [18:0] Wgt_0_555, // sfix19_En18 
  input [18:0] Wgt_0_556, // sfix19_En18 
  input [18:0] Wgt_0_557, // sfix19_En18 
  input [18:0] Wgt_0_558, // sfix19_En18 
  input [18:0] Wgt_0_559, // sfix19_En18 
  input [18:0] Wgt_0_560, // sfix19_En18 
  input [18:0] Wgt_0_561, // sfix19_En18 
  input [18:0] Wgt_0_562, // sfix19_En18 
  input [18:0] Wgt_0_563, // sfix19_En18 
  input [18:0] Wgt_0_564, // sfix19_En18 
  input [18:0] Wgt_0_565, // sfix19_En18 
  input [18:0] Wgt_0_566, // sfix19_En18 
  input [18:0] Wgt_0_567, // sfix19_En18 
  input [18:0] Wgt_0_568, // sfix19_En18 
  input [18:0] Wgt_0_569, // sfix19_En18 
  input [18:0] Wgt_0_570, // sfix19_En18 
  input [18:0] Wgt_0_571, // sfix19_En18 
  input [18:0] Wgt_0_572, // sfix19_En18 
  input [18:0] Wgt_0_573, // sfix19_En18 
  input [18:0] Wgt_0_574, // sfix19_En18 
  input [18:0] Wgt_0_575, // sfix19_En18 
  input [18:0] Wgt_0_576, // sfix19_En18 
  input [18:0] Wgt_0_577, // sfix19_En18 
  input [18:0] Wgt_0_578, // sfix19_En18 
  input [18:0] Wgt_0_579, // sfix19_En18 
  input [18:0] Wgt_0_580, // sfix19_En18 
  input [18:0] Wgt_0_581, // sfix19_En18 
  input [18:0] Wgt_0_582, // sfix19_En18 
  input [18:0] Wgt_0_583, // sfix19_En18 
  input [18:0] Wgt_0_584, // sfix19_En18 
  input [18:0] Wgt_0_585, // sfix19_En18 
  input [18:0] Wgt_0_586, // sfix19_En18 
  input [18:0] Wgt_0_587, // sfix19_En18 
  input [18:0] Wgt_0_588, // sfix19_En18 
  input [18:0] Wgt_0_589, // sfix19_En18 
  input [18:0] Wgt_0_590, // sfix19_En18 
  input [18:0] Wgt_0_591, // sfix19_En18 
  input [18:0] Wgt_0_592, // sfix19_En18 
  input [18:0] Wgt_0_593, // sfix19_En18 
  input [18:0] Wgt_0_594, // sfix19_En18 
  input [18:0] Wgt_0_595, // sfix19_En18 
  input [18:0] Wgt_0_596, // sfix19_En18 
  input [18:0] Wgt_0_597, // sfix19_En18 
  input [18:0] Wgt_0_598, // sfix19_En18 
  input [18:0] Wgt_0_599, // sfix19_En18 
  input [18:0] Wgt_0_600, // sfix19_En18 
  input [18:0] Wgt_0_601, // sfix19_En18 
  input [18:0] Wgt_0_602, // sfix19_En18 
  input [18:0] Wgt_0_603, // sfix19_En18 
  input [18:0] Wgt_0_604, // sfix19_En18 
  input [18:0] Wgt_0_605, // sfix19_En18 
  input [18:0] Wgt_0_606, // sfix19_En18 
  input [18:0] Wgt_0_607, // sfix19_En18 
  input [18:0] Wgt_0_608, // sfix19_En18 
  input [18:0] Wgt_0_609, // sfix19_En18 
  input [18:0] Wgt_0_610, // sfix19_En18 
  input [18:0] Wgt_0_611, // sfix19_En18 
  input [18:0] Wgt_0_612, // sfix19_En18 
  input [18:0] Wgt_0_613, // sfix19_En18 
  input [18:0] Wgt_0_614, // sfix19_En18 
  input [18:0] Wgt_0_615, // sfix19_En18 
  input [18:0] Wgt_0_616, // sfix19_En18 
  input [18:0] Wgt_0_617, // sfix19_En18 
  input [18:0] Wgt_0_618, // sfix19_En18 
  input [18:0] Wgt_0_619, // sfix19_En18 
  input [18:0] Wgt_0_620, // sfix19_En18 
  input [18:0] Wgt_0_621, // sfix19_En18 
  input [18:0] Wgt_0_622, // sfix19_En18 
  input [18:0] Wgt_0_623, // sfix19_En18 
  input [18:0] Wgt_0_624, // sfix19_En18 
  input [18:0] Wgt_0_625, // sfix19_En18 
  input [18:0] Wgt_0_626, // sfix19_En18 
  input [18:0] Wgt_0_627, // sfix19_En18 
  input [18:0] Wgt_0_628, // sfix19_En18 
  input [18:0] Wgt_0_629, // sfix19_En18 
  input [18:0] Wgt_0_630, // sfix19_En18 
  input [18:0] Wgt_0_631, // sfix19_En18 
  input [18:0] Wgt_0_632, // sfix19_En18 
  input [18:0] Wgt_0_633, // sfix19_En18 
  input [18:0] Wgt_0_634, // sfix19_En18 
  input [18:0] Wgt_0_635, // sfix19_En18 
  input [18:0] Wgt_0_636, // sfix19_En18 
  input [18:0] Wgt_0_637, // sfix19_En18 
  input [18:0] Wgt_0_638, // sfix19_En18 
  input [18:0] Wgt_0_639, // sfix19_En18 
  input [18:0] Wgt_0_640, // sfix19_En18 
  input [18:0] Wgt_0_641, // sfix19_En18 
  input [18:0] Wgt_0_642, // sfix19_En18 
  input [18:0] Wgt_0_643, // sfix19_En18 
  input [18:0] Wgt_0_644, // sfix19_En18 
  input [18:0] Wgt_0_645, // sfix19_En18 
  input [18:0] Wgt_0_646, // sfix19_En18 
  input [18:0] Wgt_0_647, // sfix19_En18 
  input [18:0] Wgt_0_648, // sfix19_En18 
  input [18:0] Wgt_0_649, // sfix19_En18 
  input [18:0] Wgt_0_650, // sfix19_En18 
  input [18:0] Wgt_0_651, // sfix19_En18 
  input [18:0] Wgt_0_652, // sfix19_En18 
  input [18:0] Wgt_0_653, // sfix19_En18 
  input [18:0] Wgt_0_654, // sfix19_En18 
  input [18:0] Wgt_0_655, // sfix19_En18 
  input [18:0] Wgt_0_656, // sfix19_En18 
  input [18:0] Wgt_0_657, // sfix19_En18 
  input [18:0] Wgt_0_658, // sfix19_En18 
  input [18:0] Wgt_0_659, // sfix19_En18 
  input [18:0] Wgt_0_660, // sfix19_En18 
  input [18:0] Wgt_0_661, // sfix19_En18 
  input [18:0] Wgt_0_662, // sfix19_En18 
  input [18:0] Wgt_0_663, // sfix19_En18 
  input [18:0] Wgt_0_664, // sfix19_En18 
  input [18:0] Wgt_0_665, // sfix19_En18 
  input [18:0] Wgt_0_666, // sfix19_En18 
  input [18:0] Wgt_0_667, // sfix19_En18 
  input [18:0] Wgt_0_668, // sfix19_En18 
  input [18:0] Wgt_0_669, // sfix19_En18 
  input [18:0] Wgt_0_670, // sfix19_En18 
  input [18:0] Wgt_0_671, // sfix19_En18 
  input [18:0] Wgt_0_672, // sfix19_En18 
  input [18:0] Wgt_0_673, // sfix19_En18 
  input [18:0] Wgt_0_674, // sfix19_En18 
  input [18:0] Wgt_0_675, // sfix19_En18 
  input [18:0] Wgt_0_676, // sfix19_En18 
  input [18:0] Wgt_0_677, // sfix19_En18 
  input [18:0] Wgt_0_678, // sfix19_En18 
  input [18:0] Wgt_0_679, // sfix19_En18 
  input [18:0] Wgt_0_680, // sfix19_En18 
  input [18:0] Wgt_0_681, // sfix19_En18 
  input [18:0] Wgt_0_682, // sfix19_En18 
  input [18:0] Wgt_0_683, // sfix19_En18 
  input [18:0] Wgt_0_684, // sfix19_En18 
  input [18:0] Wgt_0_685, // sfix19_En18 
  input [18:0] Wgt_0_686, // sfix19_En18 
  input [18:0] Wgt_0_687, // sfix19_En18 
  input [18:0] Wgt_0_688, // sfix19_En18 
  input [18:0] Wgt_0_689, // sfix19_En18 
  input [18:0] Wgt_0_690, // sfix19_En18 
  input [18:0] Wgt_0_691, // sfix19_En18 
  input [18:0] Wgt_0_692, // sfix19_En18 
  input [18:0] Wgt_0_693, // sfix19_En18 
  input [18:0] Wgt_0_694, // sfix19_En18 
  input [18:0] Wgt_0_695, // sfix19_En18 
  input [18:0] Wgt_0_696, // sfix19_En18 
  input [18:0] Wgt_0_697, // sfix19_En18 
  input [18:0] Wgt_0_698, // sfix19_En18 
  input [18:0] Wgt_0_699, // sfix19_En18 
  input [18:0] Wgt_0_700, // sfix19_En18 
  input [18:0] Wgt_0_701, // sfix19_En18 
  input [18:0] Wgt_0_702, // sfix19_En18 
  input [18:0] Wgt_0_703, // sfix19_En18 
  input [18:0] Wgt_0_704, // sfix19_En18 
  input [18:0] Wgt_0_705, // sfix19_En18 
  input [18:0] Wgt_0_706, // sfix19_En18 
  input [18:0] Wgt_0_707, // sfix19_En18 
  input [18:0] Wgt_0_708, // sfix19_En18 
  input [18:0] Wgt_0_709, // sfix19_En18 
  input [18:0] Wgt_0_710, // sfix19_En18 
  input [18:0] Wgt_0_711, // sfix19_En18 
  input [18:0] Wgt_0_712, // sfix19_En18 
  input [18:0] Wgt_0_713, // sfix19_En18 
  input [18:0] Wgt_0_714, // sfix19_En18 
  input [18:0] Wgt_0_715, // sfix19_En18 
  input [18:0] Wgt_0_716, // sfix19_En18 
  input [18:0] Wgt_0_717, // sfix19_En18 
  input [18:0] Wgt_0_718, // sfix19_En18 
  input [18:0] Wgt_0_719, // sfix19_En18 
  input [18:0] Wgt_0_720, // sfix19_En18 
  input [18:0] Wgt_0_721, // sfix19_En18 
  input [18:0] Wgt_0_722, // sfix19_En18 
  input [18:0] Wgt_0_723, // sfix19_En18 
  input [18:0] Wgt_0_724, // sfix19_En18 
  input [18:0] Wgt_0_725, // sfix19_En18 
  input [18:0] Wgt_0_726, // sfix19_En18 
  input [18:0] Wgt_0_727, // sfix19_En18 
  input [18:0] Wgt_0_728, // sfix19_En18 
  input [18:0] Wgt_0_729, // sfix19_En18 
  input [18:0] Wgt_0_730, // sfix19_En18 
  input [18:0] Wgt_0_731, // sfix19_En18 
  input [18:0] Wgt_0_732, // sfix19_En18 
  input [18:0] Wgt_0_733, // sfix19_En18 
  input [18:0] Wgt_0_734, // sfix19_En18 
  input [18:0] Wgt_0_735, // sfix19_En18 
  input [18:0] Wgt_0_736, // sfix19_En18 
  input [18:0] Wgt_0_737, // sfix19_En18 
  input [18:0] Wgt_0_738, // sfix19_En18 
  input [18:0] Wgt_0_739, // sfix19_En18 
  input [18:0] Wgt_0_740, // sfix19_En18 
  input [18:0] Wgt_0_741, // sfix19_En18 
  input [18:0] Wgt_0_742, // sfix19_En18 
  input [18:0] Wgt_0_743, // sfix19_En18 
  input [18:0] Wgt_0_744, // sfix19_En18 
  input [18:0] Wgt_0_745, // sfix19_En18 
  input [18:0] Wgt_0_746, // sfix19_En18 
  input [18:0] Wgt_0_747, // sfix19_En18 
  input [18:0] Wgt_0_748, // sfix19_En18 
  input [18:0] Wgt_0_749, // sfix19_En18 
  input [18:0] Wgt_0_750, // sfix19_En18 
  input [18:0] Wgt_0_751, // sfix19_En18 
  input [18:0] Wgt_0_752, // sfix19_En18 
  input [18:0] Wgt_0_753, // sfix19_En18 
  input [18:0] Wgt_0_754, // sfix19_En18 
  input [18:0] Wgt_0_755, // sfix19_En18 
  input [18:0] Wgt_0_756, // sfix19_En18 
  input [18:0] Wgt_0_757, // sfix19_En18 
  input [18:0] Wgt_0_758, // sfix19_En18 
  input [18:0] Wgt_0_759, // sfix19_En18 
  input [18:0] Wgt_0_760, // sfix19_En18 
  input [18:0] Wgt_0_761, // sfix19_En18 
  input [18:0] Wgt_0_762, // sfix19_En18 
  input [18:0] Wgt_0_763, // sfix19_En18 
  input [18:0] Wgt_0_764, // sfix19_En18 
  input [18:0] Wgt_0_765, // sfix19_En18 
  input [18:0] Wgt_0_766, // sfix19_En18 
  input [18:0] Wgt_0_767, // sfix19_En18 
  input [18:0] Wgt_0_768, // sfix19_En18 
  input [18:0] Wgt_0_769, // sfix19_En18 
  input [18:0] Wgt_0_770, // sfix19_En18 
  input [18:0] Wgt_0_771, // sfix19_En18 
  input [18:0] Wgt_0_772, // sfix19_En18 
  input [18:0] Wgt_0_773, // sfix19_En18 
  input [18:0] Wgt_0_774, // sfix19_En18 
  input [18:0] Wgt_0_775, // sfix19_En18 
  input [18:0] Wgt_0_776, // sfix19_En18 
  input [18:0] Wgt_0_777, // sfix19_En18 
  input [18:0] Wgt_0_778, // sfix19_En18 
  input [18:0] Wgt_0_779, // sfix19_En18 
  input [18:0] Wgt_0_780, // sfix19_En18 
  input [18:0] Wgt_0_781, // sfix19_En18 
  input [18:0] Wgt_0_782, // sfix19_En18 
  input [18:0] Wgt_0_783, // sfix19_En18 
  input [18:0] Wgt_0_784, // sfix19_En18 
  input [18:0] Wgt_1_0, // sfix19_En18 
  input [18:0] Wgt_1_1, // sfix19_En18 
  input [18:0] Wgt_1_2, // sfix19_En18 
  input [18:0] Wgt_1_3, // sfix19_En18 
  input [18:0] Wgt_1_4, // sfix19_En18 
  input [18:0] Wgt_1_5, // sfix19_En18 
  input [18:0] Wgt_1_6, // sfix19_En18 
  input [18:0] Wgt_1_7, // sfix19_En18 
  input [18:0] Wgt_1_8, // sfix19_En18 
  input [18:0] Wgt_1_9, // sfix19_En18 
  input [18:0] Wgt_1_10, // sfix19_En18 
  input [18:0] Wgt_1_11, // sfix19_En18 
  input [18:0] Wgt_1_12, // sfix19_En18 
  input [18:0] Wgt_1_13, // sfix19_En18 
  input [18:0] Wgt_1_14, // sfix19_En18 
  input [18:0] Wgt_1_15, // sfix19_En18 
  input [18:0] Wgt_1_16, // sfix19_En18 
  input [18:0] Wgt_1_17, // sfix19_En18 
  input [18:0] Wgt_1_18, // sfix19_En18 
  input [18:0] Wgt_1_19, // sfix19_En18 
  input [18:0] Wgt_1_20, // sfix19_En18 
  input [18:0] Wgt_1_21, // sfix19_En18 
  input [18:0] Wgt_1_22, // sfix19_En18 
  input [18:0] Wgt_1_23, // sfix19_En18 
  input [18:0] Wgt_1_24, // sfix19_En18 
  input [18:0] Wgt_1_25, // sfix19_En18 
  input [18:0] Wgt_1_26, // sfix19_En18 
  input [18:0] Wgt_1_27, // sfix19_En18 
  input [18:0] Wgt_1_28, // sfix19_En18 
  input [18:0] Wgt_1_29, // sfix19_En18 
  input [18:0] Wgt_1_30, // sfix19_En18 
  input [18:0] Wgt_1_31, // sfix19_En18 
  input [18:0] Wgt_1_32, // sfix19_En18 
  input [18:0] Wgt_1_33, // sfix19_En18 
  input [18:0] Wgt_1_34, // sfix19_En18 
  input [18:0] Wgt_1_35, // sfix19_En18 
  input [18:0] Wgt_1_36, // sfix19_En18 
  input [18:0] Wgt_1_37, // sfix19_En18 
  input [18:0] Wgt_1_38, // sfix19_En18 
  input [18:0] Wgt_1_39, // sfix19_En18 
  input [18:0] Wgt_1_40, // sfix19_En18 
  input [18:0] Wgt_1_41, // sfix19_En18 
  input [18:0] Wgt_1_42, // sfix19_En18 
  input [18:0] Wgt_1_43, // sfix19_En18 
  input [18:0] Wgt_1_44, // sfix19_En18 
  input [18:0] Wgt_1_45, // sfix19_En18 
  input [18:0] Wgt_1_46, // sfix19_En18 
  input [18:0] Wgt_1_47, // sfix19_En18 
  input [18:0] Wgt_1_48, // sfix19_En18 
  input [18:0] Wgt_1_49, // sfix19_En18 
  input [18:0] Wgt_1_50, // sfix19_En18 
  input [18:0] Wgt_1_51, // sfix19_En18 
  input [18:0] Wgt_1_52, // sfix19_En18 
  input [18:0] Wgt_1_53, // sfix19_En18 
  input [18:0] Wgt_1_54, // sfix19_En18 
  input [18:0] Wgt_1_55, // sfix19_En18 
  input [18:0] Wgt_1_56, // sfix19_En18 
  input [18:0] Wgt_1_57, // sfix19_En18 
  input [18:0] Wgt_1_58, // sfix19_En18 
  input [18:0] Wgt_1_59, // sfix19_En18 
  input [18:0] Wgt_1_60, // sfix19_En18 
  input [18:0] Wgt_1_61, // sfix19_En18 
  input [18:0] Wgt_1_62, // sfix19_En18 
  input [18:0] Wgt_1_63, // sfix19_En18 
  input [18:0] Wgt_1_64, // sfix19_En18 
  input [18:0] Wgt_1_65, // sfix19_En18 
  input [18:0] Wgt_1_66, // sfix19_En18 
  input [18:0] Wgt_1_67, // sfix19_En18 
  input [18:0] Wgt_1_68, // sfix19_En18 
  input [18:0] Wgt_1_69, // sfix19_En18 
  input [18:0] Wgt_1_70, // sfix19_En18 
  input [18:0] Wgt_1_71, // sfix19_En18 
  input [18:0] Wgt_1_72, // sfix19_En18 
  input [18:0] Wgt_1_73, // sfix19_En18 
  input [18:0] Wgt_1_74, // sfix19_En18 
  input [18:0] Wgt_1_75, // sfix19_En18 
  input [18:0] Wgt_1_76, // sfix19_En18 
  input [18:0] Wgt_1_77, // sfix19_En18 
  input [18:0] Wgt_1_78, // sfix19_En18 
  input [18:0] Wgt_1_79, // sfix19_En18 
  input [18:0] Wgt_1_80, // sfix19_En18 
  input [18:0] Wgt_1_81, // sfix19_En18 
  input [18:0] Wgt_1_82, // sfix19_En18 
  input [18:0] Wgt_1_83, // sfix19_En18 
  input [18:0] Wgt_1_84, // sfix19_En18 
  input [18:0] Wgt_1_85, // sfix19_En18 
  input [18:0] Wgt_1_86, // sfix19_En18 
  input [18:0] Wgt_1_87, // sfix19_En18 
  input [18:0] Wgt_1_88, // sfix19_En18 
  input [18:0] Wgt_1_89, // sfix19_En18 
  input [18:0] Wgt_1_90, // sfix19_En18 
  input [18:0] Wgt_1_91, // sfix19_En18 
  input [18:0] Wgt_1_92, // sfix19_En18 
  input [18:0] Wgt_1_93, // sfix19_En18 
  input [18:0] Wgt_1_94, // sfix19_En18 
  input [18:0] Wgt_1_95, // sfix19_En18 
  input [18:0] Wgt_1_96, // sfix19_En18 
  input [18:0] Wgt_1_97, // sfix19_En18 
  input [18:0] Wgt_1_98, // sfix19_En18 
  input [18:0] Wgt_1_99, // sfix19_En18 
  input [18:0] Wgt_1_100, // sfix19_En18 
  input [18:0] Wgt_1_101, // sfix19_En18 
  input [18:0] Wgt_1_102, // sfix19_En18 
  input [18:0] Wgt_1_103, // sfix19_En18 
  input [18:0] Wgt_1_104, // sfix19_En18 
  input [18:0] Wgt_1_105, // sfix19_En18 
  input [18:0] Wgt_1_106, // sfix19_En18 
  input [18:0] Wgt_1_107, // sfix19_En18 
  input [18:0] Wgt_1_108, // sfix19_En18 
  input [18:0] Wgt_1_109, // sfix19_En18 
  input [18:0] Wgt_1_110, // sfix19_En18 
  input [18:0] Wgt_1_111, // sfix19_En18 
  input [18:0] Wgt_1_112, // sfix19_En18 
  input [18:0] Wgt_1_113, // sfix19_En18 
  input [18:0] Wgt_1_114, // sfix19_En18 
  input [18:0] Wgt_1_115, // sfix19_En18 
  input [18:0] Wgt_1_116, // sfix19_En18 
  input [18:0] Wgt_1_117, // sfix19_En18 
  input [18:0] Wgt_1_118, // sfix19_En18 
  input [18:0] Wgt_1_119, // sfix19_En18 
  input [18:0] Wgt_1_120, // sfix19_En18 
  input [18:0] Wgt_1_121, // sfix19_En18 
  input [18:0] Wgt_1_122, // sfix19_En18 
  input [18:0] Wgt_1_123, // sfix19_En18 
  input [18:0] Wgt_1_124, // sfix19_En18 
  input [18:0] Wgt_1_125, // sfix19_En18 
  input [18:0] Wgt_1_126, // sfix19_En18 
  input [18:0] Wgt_1_127, // sfix19_En18 
  input [18:0] Wgt_1_128, // sfix19_En18 
  input [18:0] Wgt_1_129, // sfix19_En18 
  input [18:0] Wgt_1_130, // sfix19_En18 
  input [18:0] Wgt_1_131, // sfix19_En18 
  input [18:0] Wgt_1_132, // sfix19_En18 
  input [18:0] Wgt_1_133, // sfix19_En18 
  input [18:0] Wgt_1_134, // sfix19_En18 
  input [18:0] Wgt_1_135, // sfix19_En18 
  input [18:0] Wgt_1_136, // sfix19_En18 
  input [18:0] Wgt_1_137, // sfix19_En18 
  input [18:0] Wgt_1_138, // sfix19_En18 
  input [18:0] Wgt_1_139, // sfix19_En18 
  input [18:0] Wgt_1_140, // sfix19_En18 
  input [18:0] Wgt_1_141, // sfix19_En18 
  input [18:0] Wgt_1_142, // sfix19_En18 
  input [18:0] Wgt_1_143, // sfix19_En18 
  input [18:0] Wgt_1_144, // sfix19_En18 
  input [18:0] Wgt_1_145, // sfix19_En18 
  input [18:0] Wgt_1_146, // sfix19_En18 
  input [18:0] Wgt_1_147, // sfix19_En18 
  input [18:0] Wgt_1_148, // sfix19_En18 
  input [18:0] Wgt_1_149, // sfix19_En18 
  input [18:0] Wgt_1_150, // sfix19_En18 
  input [18:0] Wgt_1_151, // sfix19_En18 
  input [18:0] Wgt_1_152, // sfix19_En18 
  input [18:0] Wgt_1_153, // sfix19_En18 
  input [18:0] Wgt_1_154, // sfix19_En18 
  input [18:0] Wgt_1_155, // sfix19_En18 
  input [18:0] Wgt_1_156, // sfix19_En18 
  input [18:0] Wgt_1_157, // sfix19_En18 
  input [18:0] Wgt_1_158, // sfix19_En18 
  input [18:0] Wgt_1_159, // sfix19_En18 
  input [18:0] Wgt_1_160, // sfix19_En18 
  input [18:0] Wgt_1_161, // sfix19_En18 
  input [18:0] Wgt_1_162, // sfix19_En18 
  input [18:0] Wgt_1_163, // sfix19_En18 
  input [18:0] Wgt_1_164, // sfix19_En18 
  input [18:0] Wgt_1_165, // sfix19_En18 
  input [18:0] Wgt_1_166, // sfix19_En18 
  input [18:0] Wgt_1_167, // sfix19_En18 
  input [18:0] Wgt_1_168, // sfix19_En18 
  input [18:0] Wgt_1_169, // sfix19_En18 
  input [18:0] Wgt_1_170, // sfix19_En18 
  input [18:0] Wgt_1_171, // sfix19_En18 
  input [18:0] Wgt_1_172, // sfix19_En18 
  input [18:0] Wgt_1_173, // sfix19_En18 
  input [18:0] Wgt_1_174, // sfix19_En18 
  input [18:0] Wgt_1_175, // sfix19_En18 
  input [18:0] Wgt_1_176, // sfix19_En18 
  input [18:0] Wgt_1_177, // sfix19_En18 
  input [18:0] Wgt_1_178, // sfix19_En18 
  input [18:0] Wgt_1_179, // sfix19_En18 
  input [18:0] Wgt_1_180, // sfix19_En18 
  input [18:0] Wgt_1_181, // sfix19_En18 
  input [18:0] Wgt_1_182, // sfix19_En18 
  input [18:0] Wgt_1_183, // sfix19_En18 
  input [18:0] Wgt_1_184, // sfix19_En18 
  input [18:0] Wgt_1_185, // sfix19_En18 
  input [18:0] Wgt_1_186, // sfix19_En18 
  input [18:0] Wgt_1_187, // sfix19_En18 
  input [18:0] Wgt_1_188, // sfix19_En18 
  input [18:0] Wgt_1_189, // sfix19_En18 
  input [18:0] Wgt_1_190, // sfix19_En18 
  input [18:0] Wgt_1_191, // sfix19_En18 
  input [18:0] Wgt_1_192, // sfix19_En18 
  input [18:0] Wgt_1_193, // sfix19_En18 
  input [18:0] Wgt_1_194, // sfix19_En18 
  input [18:0] Wgt_1_195, // sfix19_En18 
  input [18:0] Wgt_1_196, // sfix19_En18 
  input [18:0] Wgt_1_197, // sfix19_En18 
  input [18:0] Wgt_1_198, // sfix19_En18 
  input [18:0] Wgt_1_199, // sfix19_En18 
  input [18:0] Wgt_1_200, // sfix19_En18 
  input [18:0] Wgt_1_201, // sfix19_En18 
  input [18:0] Wgt_1_202, // sfix19_En18 
  input [18:0] Wgt_1_203, // sfix19_En18 
  input [18:0] Wgt_1_204, // sfix19_En18 
  input [18:0] Wgt_1_205, // sfix19_En18 
  input [18:0] Wgt_1_206, // sfix19_En18 
  input [18:0] Wgt_1_207, // sfix19_En18 
  input [18:0] Wgt_1_208, // sfix19_En18 
  input [18:0] Wgt_1_209, // sfix19_En18 
  input [18:0] Wgt_1_210, // sfix19_En18 
  input [18:0] Wgt_1_211, // sfix19_En18 
  input [18:0] Wgt_1_212, // sfix19_En18 
  input [18:0] Wgt_1_213, // sfix19_En18 
  input [18:0] Wgt_1_214, // sfix19_En18 
  input [18:0] Wgt_1_215, // sfix19_En18 
  input [18:0] Wgt_1_216, // sfix19_En18 
  input [18:0] Wgt_1_217, // sfix19_En18 
  input [18:0] Wgt_1_218, // sfix19_En18 
  input [18:0] Wgt_1_219, // sfix19_En18 
  input [18:0] Wgt_1_220, // sfix19_En18 
  input [18:0] Wgt_1_221, // sfix19_En18 
  input [18:0] Wgt_1_222, // sfix19_En18 
  input [18:0] Wgt_1_223, // sfix19_En18 
  input [18:0] Wgt_1_224, // sfix19_En18 
  input [18:0] Wgt_1_225, // sfix19_En18 
  input [18:0] Wgt_1_226, // sfix19_En18 
  input [18:0] Wgt_1_227, // sfix19_En18 
  input [18:0] Wgt_1_228, // sfix19_En18 
  input [18:0] Wgt_1_229, // sfix19_En18 
  input [18:0] Wgt_1_230, // sfix19_En18 
  input [18:0] Wgt_1_231, // sfix19_En18 
  input [18:0] Wgt_1_232, // sfix19_En18 
  input [18:0] Wgt_1_233, // sfix19_En18 
  input [18:0] Wgt_1_234, // sfix19_En18 
  input [18:0] Wgt_1_235, // sfix19_En18 
  input [18:0] Wgt_1_236, // sfix19_En18 
  input [18:0] Wgt_1_237, // sfix19_En18 
  input [18:0] Wgt_1_238, // sfix19_En18 
  input [18:0] Wgt_1_239, // sfix19_En18 
  input [18:0] Wgt_1_240, // sfix19_En18 
  input [18:0] Wgt_1_241, // sfix19_En18 
  input [18:0] Wgt_1_242, // sfix19_En18 
  input [18:0] Wgt_1_243, // sfix19_En18 
  input [18:0] Wgt_1_244, // sfix19_En18 
  input [18:0] Wgt_1_245, // sfix19_En18 
  input [18:0] Wgt_1_246, // sfix19_En18 
  input [18:0] Wgt_1_247, // sfix19_En18 
  input [18:0] Wgt_1_248, // sfix19_En18 
  input [18:0] Wgt_1_249, // sfix19_En18 
  input [18:0] Wgt_1_250, // sfix19_En18 
  input [18:0] Wgt_1_251, // sfix19_En18 
  input [18:0] Wgt_1_252, // sfix19_En18 
  input [18:0] Wgt_1_253, // sfix19_En18 
  input [18:0] Wgt_1_254, // sfix19_En18 
  input [18:0] Wgt_1_255, // sfix19_En18 
  input [18:0] Wgt_1_256, // sfix19_En18 
  input [18:0] Wgt_1_257, // sfix19_En18 
  input [18:0] Wgt_1_258, // sfix19_En18 
  input [18:0] Wgt_1_259, // sfix19_En18 
  input [18:0] Wgt_1_260, // sfix19_En18 
  input [18:0] Wgt_1_261, // sfix19_En18 
  input [18:0] Wgt_1_262, // sfix19_En18 
  input [18:0] Wgt_1_263, // sfix19_En18 
  input [18:0] Wgt_1_264, // sfix19_En18 
  input [18:0] Wgt_1_265, // sfix19_En18 
  input [18:0] Wgt_1_266, // sfix19_En18 
  input [18:0] Wgt_1_267, // sfix19_En18 
  input [18:0] Wgt_1_268, // sfix19_En18 
  input [18:0] Wgt_1_269, // sfix19_En18 
  input [18:0] Wgt_1_270, // sfix19_En18 
  input [18:0] Wgt_1_271, // sfix19_En18 
  input [18:0] Wgt_1_272, // sfix19_En18 
  input [18:0] Wgt_1_273, // sfix19_En18 
  input [18:0] Wgt_1_274, // sfix19_En18 
  input [18:0] Wgt_1_275, // sfix19_En18 
  input [18:0] Wgt_1_276, // sfix19_En18 
  input [18:0] Wgt_1_277, // sfix19_En18 
  input [18:0] Wgt_1_278, // sfix19_En18 
  input [18:0] Wgt_1_279, // sfix19_En18 
  input [18:0] Wgt_1_280, // sfix19_En18 
  input [18:0] Wgt_1_281, // sfix19_En18 
  input [18:0] Wgt_1_282, // sfix19_En18 
  input [18:0] Wgt_1_283, // sfix19_En18 
  input [18:0] Wgt_1_284, // sfix19_En18 
  input [18:0] Wgt_1_285, // sfix19_En18 
  input [18:0] Wgt_1_286, // sfix19_En18 
  input [18:0] Wgt_1_287, // sfix19_En18 
  input [18:0] Wgt_1_288, // sfix19_En18 
  input [18:0] Wgt_1_289, // sfix19_En18 
  input [18:0] Wgt_1_290, // sfix19_En18 
  input [18:0] Wgt_1_291, // sfix19_En18 
  input [18:0] Wgt_1_292, // sfix19_En18 
  input [18:0] Wgt_1_293, // sfix19_En18 
  input [18:0] Wgt_1_294, // sfix19_En18 
  input [18:0] Wgt_1_295, // sfix19_En18 
  input [18:0] Wgt_1_296, // sfix19_En18 
  input [18:0] Wgt_1_297, // sfix19_En18 
  input [18:0] Wgt_1_298, // sfix19_En18 
  input [18:0] Wgt_1_299, // sfix19_En18 
  input [18:0] Wgt_1_300, // sfix19_En18 
  input [18:0] Wgt_1_301, // sfix19_En18 
  input [18:0] Wgt_1_302, // sfix19_En18 
  input [18:0] Wgt_1_303, // sfix19_En18 
  input [18:0] Wgt_1_304, // sfix19_En18 
  input [18:0] Wgt_1_305, // sfix19_En18 
  input [18:0] Wgt_1_306, // sfix19_En18 
  input [18:0] Wgt_1_307, // sfix19_En18 
  input [18:0] Wgt_1_308, // sfix19_En18 
  input [18:0] Wgt_1_309, // sfix19_En18 
  input [18:0] Wgt_1_310, // sfix19_En18 
  input [18:0] Wgt_1_311, // sfix19_En18 
  input [18:0] Wgt_1_312, // sfix19_En18 
  input [18:0] Wgt_1_313, // sfix19_En18 
  input [18:0] Wgt_1_314, // sfix19_En18 
  input [18:0] Wgt_1_315, // sfix19_En18 
  input [18:0] Wgt_1_316, // sfix19_En18 
  input [18:0] Wgt_1_317, // sfix19_En18 
  input [18:0] Wgt_1_318, // sfix19_En18 
  input [18:0] Wgt_1_319, // sfix19_En18 
  input [18:0] Wgt_1_320, // sfix19_En18 
  input [18:0] Wgt_1_321, // sfix19_En18 
  input [18:0] Wgt_1_322, // sfix19_En18 
  input [18:0] Wgt_1_323, // sfix19_En18 
  input [18:0] Wgt_1_324, // sfix19_En18 
  input [18:0] Wgt_1_325, // sfix19_En18 
  input [18:0] Wgt_1_326, // sfix19_En18 
  input [18:0] Wgt_1_327, // sfix19_En18 
  input [18:0] Wgt_1_328, // sfix19_En18 
  input [18:0] Wgt_1_329, // sfix19_En18 
  input [18:0] Wgt_1_330, // sfix19_En18 
  input [18:0] Wgt_1_331, // sfix19_En18 
  input [18:0] Wgt_1_332, // sfix19_En18 
  input [18:0] Wgt_1_333, // sfix19_En18 
  input [18:0] Wgt_1_334, // sfix19_En18 
  input [18:0] Wgt_1_335, // sfix19_En18 
  input [18:0] Wgt_1_336, // sfix19_En18 
  input [18:0] Wgt_1_337, // sfix19_En18 
  input [18:0] Wgt_1_338, // sfix19_En18 
  input [18:0] Wgt_1_339, // sfix19_En18 
  input [18:0] Wgt_1_340, // sfix19_En18 
  input [18:0] Wgt_1_341, // sfix19_En18 
  input [18:0] Wgt_1_342, // sfix19_En18 
  input [18:0] Wgt_1_343, // sfix19_En18 
  input [18:0] Wgt_1_344, // sfix19_En18 
  input [18:0] Wgt_1_345, // sfix19_En18 
  input [18:0] Wgt_1_346, // sfix19_En18 
  input [18:0] Wgt_1_347, // sfix19_En18 
  input [18:0] Wgt_1_348, // sfix19_En18 
  input [18:0] Wgt_1_349, // sfix19_En18 
  input [18:0] Wgt_1_350, // sfix19_En18 
  input [18:0] Wgt_1_351, // sfix19_En18 
  input [18:0] Wgt_1_352, // sfix19_En18 
  input [18:0] Wgt_1_353, // sfix19_En18 
  input [18:0] Wgt_1_354, // sfix19_En18 
  input [18:0] Wgt_1_355, // sfix19_En18 
  input [18:0] Wgt_1_356, // sfix19_En18 
  input [18:0] Wgt_1_357, // sfix19_En18 
  input [18:0] Wgt_1_358, // sfix19_En18 
  input [18:0] Wgt_1_359, // sfix19_En18 
  input [18:0] Wgt_1_360, // sfix19_En18 
  input [18:0] Wgt_1_361, // sfix19_En18 
  input [18:0] Wgt_1_362, // sfix19_En18 
  input [18:0] Wgt_1_363, // sfix19_En18 
  input [18:0] Wgt_1_364, // sfix19_En18 
  input [18:0] Wgt_1_365, // sfix19_En18 
  input [18:0] Wgt_1_366, // sfix19_En18 
  input [18:0] Wgt_1_367, // sfix19_En18 
  input [18:0] Wgt_1_368, // sfix19_En18 
  input [18:0] Wgt_1_369, // sfix19_En18 
  input [18:0] Wgt_1_370, // sfix19_En18 
  input [18:0] Wgt_1_371, // sfix19_En18 
  input [18:0] Wgt_1_372, // sfix19_En18 
  input [18:0] Wgt_1_373, // sfix19_En18 
  input [18:0] Wgt_1_374, // sfix19_En18 
  input [18:0] Wgt_1_375, // sfix19_En18 
  input [18:0] Wgt_1_376, // sfix19_En18 
  input [18:0] Wgt_1_377, // sfix19_En18 
  input [18:0] Wgt_1_378, // sfix19_En18 
  input [18:0] Wgt_1_379, // sfix19_En18 
  input [18:0] Wgt_1_380, // sfix19_En18 
  input [18:0] Wgt_1_381, // sfix19_En18 
  input [18:0] Wgt_1_382, // sfix19_En18 
  input [18:0] Wgt_1_383, // sfix19_En18 
  input [18:0] Wgt_1_384, // sfix19_En18 
  input [18:0] Wgt_1_385, // sfix19_En18 
  input [18:0] Wgt_1_386, // sfix19_En18 
  input [18:0] Wgt_1_387, // sfix19_En18 
  input [18:0] Wgt_1_388, // sfix19_En18 
  input [18:0] Wgt_1_389, // sfix19_En18 
  input [18:0] Wgt_1_390, // sfix19_En18 
  input [18:0] Wgt_1_391, // sfix19_En18 
  input [18:0] Wgt_1_392, // sfix19_En18 
  input [18:0] Wgt_1_393, // sfix19_En18 
  input [18:0] Wgt_1_394, // sfix19_En18 
  input [18:0] Wgt_1_395, // sfix19_En18 
  input [18:0] Wgt_1_396, // sfix19_En18 
  input [18:0] Wgt_1_397, // sfix19_En18 
  input [18:0] Wgt_1_398, // sfix19_En18 
  input [18:0] Wgt_1_399, // sfix19_En18 
  input [18:0] Wgt_1_400, // sfix19_En18 
  input [18:0] Wgt_1_401, // sfix19_En18 
  input [18:0] Wgt_1_402, // sfix19_En18 
  input [18:0] Wgt_1_403, // sfix19_En18 
  input [18:0] Wgt_1_404, // sfix19_En18 
  input [18:0] Wgt_1_405, // sfix19_En18 
  input [18:0] Wgt_1_406, // sfix19_En18 
  input [18:0] Wgt_1_407, // sfix19_En18 
  input [18:0] Wgt_1_408, // sfix19_En18 
  input [18:0] Wgt_1_409, // sfix19_En18 
  input [18:0] Wgt_1_410, // sfix19_En18 
  input [18:0] Wgt_1_411, // sfix19_En18 
  input [18:0] Wgt_1_412, // sfix19_En18 
  input [18:0] Wgt_1_413, // sfix19_En18 
  input [18:0] Wgt_1_414, // sfix19_En18 
  input [18:0] Wgt_1_415, // sfix19_En18 
  input [18:0] Wgt_1_416, // sfix19_En18 
  input [18:0] Wgt_1_417, // sfix19_En18 
  input [18:0] Wgt_1_418, // sfix19_En18 
  input [18:0] Wgt_1_419, // sfix19_En18 
  input [18:0] Wgt_1_420, // sfix19_En18 
  input [18:0] Wgt_1_421, // sfix19_En18 
  input [18:0] Wgt_1_422, // sfix19_En18 
  input [18:0] Wgt_1_423, // sfix19_En18 
  input [18:0] Wgt_1_424, // sfix19_En18 
  input [18:0] Wgt_1_425, // sfix19_En18 
  input [18:0] Wgt_1_426, // sfix19_En18 
  input [18:0] Wgt_1_427, // sfix19_En18 
  input [18:0] Wgt_1_428, // sfix19_En18 
  input [18:0] Wgt_1_429, // sfix19_En18 
  input [18:0] Wgt_1_430, // sfix19_En18 
  input [18:0] Wgt_1_431, // sfix19_En18 
  input [18:0] Wgt_1_432, // sfix19_En18 
  input [18:0] Wgt_1_433, // sfix19_En18 
  input [18:0] Wgt_1_434, // sfix19_En18 
  input [18:0] Wgt_1_435, // sfix19_En18 
  input [18:0] Wgt_1_436, // sfix19_En18 
  input [18:0] Wgt_1_437, // sfix19_En18 
  input [18:0] Wgt_1_438, // sfix19_En18 
  input [18:0] Wgt_1_439, // sfix19_En18 
  input [18:0] Wgt_1_440, // sfix19_En18 
  input [18:0] Wgt_1_441, // sfix19_En18 
  input [18:0] Wgt_1_442, // sfix19_En18 
  input [18:0] Wgt_1_443, // sfix19_En18 
  input [18:0] Wgt_1_444, // sfix19_En18 
  input [18:0] Wgt_1_445, // sfix19_En18 
  input [18:0] Wgt_1_446, // sfix19_En18 
  input [18:0] Wgt_1_447, // sfix19_En18 
  input [18:0] Wgt_1_448, // sfix19_En18 
  input [18:0] Wgt_1_449, // sfix19_En18 
  input [18:0] Wgt_1_450, // sfix19_En18 
  input [18:0] Wgt_1_451, // sfix19_En18 
  input [18:0] Wgt_1_452, // sfix19_En18 
  input [18:0] Wgt_1_453, // sfix19_En18 
  input [18:0] Wgt_1_454, // sfix19_En18 
  input [18:0] Wgt_1_455, // sfix19_En18 
  input [18:0] Wgt_1_456, // sfix19_En18 
  input [18:0] Wgt_1_457, // sfix19_En18 
  input [18:0] Wgt_1_458, // sfix19_En18 
  input [18:0] Wgt_1_459, // sfix19_En18 
  input [18:0] Wgt_1_460, // sfix19_En18 
  input [18:0] Wgt_1_461, // sfix19_En18 
  input [18:0] Wgt_1_462, // sfix19_En18 
  input [18:0] Wgt_1_463, // sfix19_En18 
  input [18:0] Wgt_1_464, // sfix19_En18 
  input [18:0] Wgt_1_465, // sfix19_En18 
  input [18:0] Wgt_1_466, // sfix19_En18 
  input [18:0] Wgt_1_467, // sfix19_En18 
  input [18:0] Wgt_1_468, // sfix19_En18 
  input [18:0] Wgt_1_469, // sfix19_En18 
  input [18:0] Wgt_1_470, // sfix19_En18 
  input [18:0] Wgt_1_471, // sfix19_En18 
  input [18:0] Wgt_1_472, // sfix19_En18 
  input [18:0] Wgt_1_473, // sfix19_En18 
  input [18:0] Wgt_1_474, // sfix19_En18 
  input [18:0] Wgt_1_475, // sfix19_En18 
  input [18:0] Wgt_1_476, // sfix19_En18 
  input [18:0] Wgt_1_477, // sfix19_En18 
  input [18:0] Wgt_1_478, // sfix19_En18 
  input [18:0] Wgt_1_479, // sfix19_En18 
  input [18:0] Wgt_1_480, // sfix19_En18 
  input [18:0] Wgt_1_481, // sfix19_En18 
  input [18:0] Wgt_1_482, // sfix19_En18 
  input [18:0] Wgt_1_483, // sfix19_En18 
  input [18:0] Wgt_1_484, // sfix19_En18 
  input [18:0] Wgt_1_485, // sfix19_En18 
  input [18:0] Wgt_1_486, // sfix19_En18 
  input [18:0] Wgt_1_487, // sfix19_En18 
  input [18:0] Wgt_1_488, // sfix19_En18 
  input [18:0] Wgt_1_489, // sfix19_En18 
  input [18:0] Wgt_1_490, // sfix19_En18 
  input [18:0] Wgt_1_491, // sfix19_En18 
  input [18:0] Wgt_1_492, // sfix19_En18 
  input [18:0] Wgt_1_493, // sfix19_En18 
  input [18:0] Wgt_1_494, // sfix19_En18 
  input [18:0] Wgt_1_495, // sfix19_En18 
  input [18:0] Wgt_1_496, // sfix19_En18 
  input [18:0] Wgt_1_497, // sfix19_En18 
  input [18:0] Wgt_1_498, // sfix19_En18 
  input [18:0] Wgt_1_499, // sfix19_En18 
  input [18:0] Wgt_1_500, // sfix19_En18 
  input [18:0] Wgt_1_501, // sfix19_En18 
  input [18:0] Wgt_1_502, // sfix19_En18 
  input [18:0] Wgt_1_503, // sfix19_En18 
  input [18:0] Wgt_1_504, // sfix19_En18 
  input [18:0] Wgt_1_505, // sfix19_En18 
  input [18:0] Wgt_1_506, // sfix19_En18 
  input [18:0] Wgt_1_507, // sfix19_En18 
  input [18:0] Wgt_1_508, // sfix19_En18 
  input [18:0] Wgt_1_509, // sfix19_En18 
  input [18:0] Wgt_1_510, // sfix19_En18 
  input [18:0] Wgt_1_511, // sfix19_En18 
  input [18:0] Wgt_1_512, // sfix19_En18 
  input [18:0] Wgt_1_513, // sfix19_En18 
  input [18:0] Wgt_1_514, // sfix19_En18 
  input [18:0] Wgt_1_515, // sfix19_En18 
  input [18:0] Wgt_1_516, // sfix19_En18 
  input [18:0] Wgt_1_517, // sfix19_En18 
  input [18:0] Wgt_1_518, // sfix19_En18 
  input [18:0] Wgt_1_519, // sfix19_En18 
  input [18:0] Wgt_1_520, // sfix19_En18 
  input [18:0] Wgt_1_521, // sfix19_En18 
  input [18:0] Wgt_1_522, // sfix19_En18 
  input [18:0] Wgt_1_523, // sfix19_En18 
  input [18:0] Wgt_1_524, // sfix19_En18 
  input [18:0] Wgt_1_525, // sfix19_En18 
  input [18:0] Wgt_1_526, // sfix19_En18 
  input [18:0] Wgt_1_527, // sfix19_En18 
  input [18:0] Wgt_1_528, // sfix19_En18 
  input [18:0] Wgt_1_529, // sfix19_En18 
  input [18:0] Wgt_1_530, // sfix19_En18 
  input [18:0] Wgt_1_531, // sfix19_En18 
  input [18:0] Wgt_1_532, // sfix19_En18 
  input [18:0] Wgt_1_533, // sfix19_En18 
  input [18:0] Wgt_1_534, // sfix19_En18 
  input [18:0] Wgt_1_535, // sfix19_En18 
  input [18:0] Wgt_1_536, // sfix19_En18 
  input [18:0] Wgt_1_537, // sfix19_En18 
  input [18:0] Wgt_1_538, // sfix19_En18 
  input [18:0] Wgt_1_539, // sfix19_En18 
  input [18:0] Wgt_1_540, // sfix19_En18 
  input [18:0] Wgt_1_541, // sfix19_En18 
  input [18:0] Wgt_1_542, // sfix19_En18 
  input [18:0] Wgt_1_543, // sfix19_En18 
  input [18:0] Wgt_1_544, // sfix19_En18 
  input [18:0] Wgt_1_545, // sfix19_En18 
  input [18:0] Wgt_1_546, // sfix19_En18 
  input [18:0] Wgt_1_547, // sfix19_En18 
  input [18:0] Wgt_1_548, // sfix19_En18 
  input [18:0] Wgt_1_549, // sfix19_En18 
  input [18:0] Wgt_1_550, // sfix19_En18 
  input [18:0] Wgt_1_551, // sfix19_En18 
  input [18:0] Wgt_1_552, // sfix19_En18 
  input [18:0] Wgt_1_553, // sfix19_En18 
  input [18:0] Wgt_1_554, // sfix19_En18 
  input [18:0] Wgt_1_555, // sfix19_En18 
  input [18:0] Wgt_1_556, // sfix19_En18 
  input [18:0] Wgt_1_557, // sfix19_En18 
  input [18:0] Wgt_1_558, // sfix19_En18 
  input [18:0] Wgt_1_559, // sfix19_En18 
  input [18:0] Wgt_1_560, // sfix19_En18 
  input [18:0] Wgt_1_561, // sfix19_En18 
  input [18:0] Wgt_1_562, // sfix19_En18 
  input [18:0] Wgt_1_563, // sfix19_En18 
  input [18:0] Wgt_1_564, // sfix19_En18 
  input [18:0] Wgt_1_565, // sfix19_En18 
  input [18:0] Wgt_1_566, // sfix19_En18 
  input [18:0] Wgt_1_567, // sfix19_En18 
  input [18:0] Wgt_1_568, // sfix19_En18 
  input [18:0] Wgt_1_569, // sfix19_En18 
  input [18:0] Wgt_1_570, // sfix19_En18 
  input [18:0] Wgt_1_571, // sfix19_En18 
  input [18:0] Wgt_1_572, // sfix19_En18 
  input [18:0] Wgt_1_573, // sfix19_En18 
  input [18:0] Wgt_1_574, // sfix19_En18 
  input [18:0] Wgt_1_575, // sfix19_En18 
  input [18:0] Wgt_1_576, // sfix19_En18 
  input [18:0] Wgt_1_577, // sfix19_En18 
  input [18:0] Wgt_1_578, // sfix19_En18 
  input [18:0] Wgt_1_579, // sfix19_En18 
  input [18:0] Wgt_1_580, // sfix19_En18 
  input [18:0] Wgt_1_581, // sfix19_En18 
  input [18:0] Wgt_1_582, // sfix19_En18 
  input [18:0] Wgt_1_583, // sfix19_En18 
  input [18:0] Wgt_1_584, // sfix19_En18 
  input [18:0] Wgt_1_585, // sfix19_En18 
  input [18:0] Wgt_1_586, // sfix19_En18 
  input [18:0] Wgt_1_587, // sfix19_En18 
  input [18:0] Wgt_1_588, // sfix19_En18 
  input [18:0] Wgt_1_589, // sfix19_En18 
  input [18:0] Wgt_1_590, // sfix19_En18 
  input [18:0] Wgt_1_591, // sfix19_En18 
  input [18:0] Wgt_1_592, // sfix19_En18 
  input [18:0] Wgt_1_593, // sfix19_En18 
  input [18:0] Wgt_1_594, // sfix19_En18 
  input [18:0] Wgt_1_595, // sfix19_En18 
  input [18:0] Wgt_1_596, // sfix19_En18 
  input [18:0] Wgt_1_597, // sfix19_En18 
  input [18:0] Wgt_1_598, // sfix19_En18 
  input [18:0] Wgt_1_599, // sfix19_En18 
  input [18:0] Wgt_1_600, // sfix19_En18 
  input [18:0] Wgt_1_601, // sfix19_En18 
  input [18:0] Wgt_1_602, // sfix19_En18 
  input [18:0] Wgt_1_603, // sfix19_En18 
  input [18:0] Wgt_1_604, // sfix19_En18 
  input [18:0] Wgt_1_605, // sfix19_En18 
  input [18:0] Wgt_1_606, // sfix19_En18 
  input [18:0] Wgt_1_607, // sfix19_En18 
  input [18:0] Wgt_1_608, // sfix19_En18 
  input [18:0] Wgt_1_609, // sfix19_En18 
  input [18:0] Wgt_1_610, // sfix19_En18 
  input [18:0] Wgt_1_611, // sfix19_En18 
  input [18:0] Wgt_1_612, // sfix19_En18 
  input [18:0] Wgt_1_613, // sfix19_En18 
  input [18:0] Wgt_1_614, // sfix19_En18 
  input [18:0] Wgt_1_615, // sfix19_En18 
  input [18:0] Wgt_1_616, // sfix19_En18 
  input [18:0] Wgt_1_617, // sfix19_En18 
  input [18:0] Wgt_1_618, // sfix19_En18 
  input [18:0] Wgt_1_619, // sfix19_En18 
  input [18:0] Wgt_1_620, // sfix19_En18 
  input [18:0] Wgt_1_621, // sfix19_En18 
  input [18:0] Wgt_1_622, // sfix19_En18 
  input [18:0] Wgt_1_623, // sfix19_En18 
  input [18:0] Wgt_1_624, // sfix19_En18 
  input [18:0] Wgt_1_625, // sfix19_En18 
  input [18:0] Wgt_1_626, // sfix19_En18 
  input [18:0] Wgt_1_627, // sfix19_En18 
  input [18:0] Wgt_1_628, // sfix19_En18 
  input [18:0] Wgt_1_629, // sfix19_En18 
  input [18:0] Wgt_1_630, // sfix19_En18 
  input [18:0] Wgt_1_631, // sfix19_En18 
  input [18:0] Wgt_1_632, // sfix19_En18 
  input [18:0] Wgt_1_633, // sfix19_En18 
  input [18:0] Wgt_1_634, // sfix19_En18 
  input [18:0] Wgt_1_635, // sfix19_En18 
  input [18:0] Wgt_1_636, // sfix19_En18 
  input [18:0] Wgt_1_637, // sfix19_En18 
  input [18:0] Wgt_1_638, // sfix19_En18 
  input [18:0] Wgt_1_639, // sfix19_En18 
  input [18:0] Wgt_1_640, // sfix19_En18 
  input [18:0] Wgt_1_641, // sfix19_En18 
  input [18:0] Wgt_1_642, // sfix19_En18 
  input [18:0] Wgt_1_643, // sfix19_En18 
  input [18:0] Wgt_1_644, // sfix19_En18 
  input [18:0] Wgt_1_645, // sfix19_En18 
  input [18:0] Wgt_1_646, // sfix19_En18 
  input [18:0] Wgt_1_647, // sfix19_En18 
  input [18:0] Wgt_1_648, // sfix19_En18 
  input [18:0] Wgt_1_649, // sfix19_En18 
  input [18:0] Wgt_1_650, // sfix19_En18 
  input [18:0] Wgt_1_651, // sfix19_En18 
  input [18:0] Wgt_1_652, // sfix19_En18 
  input [18:0] Wgt_1_653, // sfix19_En18 
  input [18:0] Wgt_1_654, // sfix19_En18 
  input [18:0] Wgt_1_655, // sfix19_En18 
  input [18:0] Wgt_1_656, // sfix19_En18 
  input [18:0] Wgt_1_657, // sfix19_En18 
  input [18:0] Wgt_1_658, // sfix19_En18 
  input [18:0] Wgt_1_659, // sfix19_En18 
  input [18:0] Wgt_1_660, // sfix19_En18 
  input [18:0] Wgt_1_661, // sfix19_En18 
  input [18:0] Wgt_1_662, // sfix19_En18 
  input [18:0] Wgt_1_663, // sfix19_En18 
  input [18:0] Wgt_1_664, // sfix19_En18 
  input [18:0] Wgt_1_665, // sfix19_En18 
  input [18:0] Wgt_1_666, // sfix19_En18 
  input [18:0] Wgt_1_667, // sfix19_En18 
  input [18:0] Wgt_1_668, // sfix19_En18 
  input [18:0] Wgt_1_669, // sfix19_En18 
  input [18:0] Wgt_1_670, // sfix19_En18 
  input [18:0] Wgt_1_671, // sfix19_En18 
  input [18:0] Wgt_1_672, // sfix19_En18 
  input [18:0] Wgt_1_673, // sfix19_En18 
  input [18:0] Wgt_1_674, // sfix19_En18 
  input [18:0] Wgt_1_675, // sfix19_En18 
  input [18:0] Wgt_1_676, // sfix19_En18 
  input [18:0] Wgt_1_677, // sfix19_En18 
  input [18:0] Wgt_1_678, // sfix19_En18 
  input [18:0] Wgt_1_679, // sfix19_En18 
  input [18:0] Wgt_1_680, // sfix19_En18 
  input [18:0] Wgt_1_681, // sfix19_En18 
  input [18:0] Wgt_1_682, // sfix19_En18 
  input [18:0] Wgt_1_683, // sfix19_En18 
  input [18:0] Wgt_1_684, // sfix19_En18 
  input [18:0] Wgt_1_685, // sfix19_En18 
  input [18:0] Wgt_1_686, // sfix19_En18 
  input [18:0] Wgt_1_687, // sfix19_En18 
  input [18:0] Wgt_1_688, // sfix19_En18 
  input [18:0] Wgt_1_689, // sfix19_En18 
  input [18:0] Wgt_1_690, // sfix19_En18 
  input [18:0] Wgt_1_691, // sfix19_En18 
  input [18:0] Wgt_1_692, // sfix19_En18 
  input [18:0] Wgt_1_693, // sfix19_En18 
  input [18:0] Wgt_1_694, // sfix19_En18 
  input [18:0] Wgt_1_695, // sfix19_En18 
  input [18:0] Wgt_1_696, // sfix19_En18 
  input [18:0] Wgt_1_697, // sfix19_En18 
  input [18:0] Wgt_1_698, // sfix19_En18 
  input [18:0] Wgt_1_699, // sfix19_En18 
  input [18:0] Wgt_1_700, // sfix19_En18 
  input [18:0] Wgt_1_701, // sfix19_En18 
  input [18:0] Wgt_1_702, // sfix19_En18 
  input [18:0] Wgt_1_703, // sfix19_En18 
  input [18:0] Wgt_1_704, // sfix19_En18 
  input [18:0] Wgt_1_705, // sfix19_En18 
  input [18:0] Wgt_1_706, // sfix19_En18 
  input [18:0] Wgt_1_707, // sfix19_En18 
  input [18:0] Wgt_1_708, // sfix19_En18 
  input [18:0] Wgt_1_709, // sfix19_En18 
  input [18:0] Wgt_1_710, // sfix19_En18 
  input [18:0] Wgt_1_711, // sfix19_En18 
  input [18:0] Wgt_1_712, // sfix19_En18 
  input [18:0] Wgt_1_713, // sfix19_En18 
  input [18:0] Wgt_1_714, // sfix19_En18 
  input [18:0] Wgt_1_715, // sfix19_En18 
  input [18:0] Wgt_1_716, // sfix19_En18 
  input [18:0] Wgt_1_717, // sfix19_En18 
  input [18:0] Wgt_1_718, // sfix19_En18 
  input [18:0] Wgt_1_719, // sfix19_En18 
  input [18:0] Wgt_1_720, // sfix19_En18 
  input [18:0] Wgt_1_721, // sfix19_En18 
  input [18:0] Wgt_1_722, // sfix19_En18 
  input [18:0] Wgt_1_723, // sfix19_En18 
  input [18:0] Wgt_1_724, // sfix19_En18 
  input [18:0] Wgt_1_725, // sfix19_En18 
  input [18:0] Wgt_1_726, // sfix19_En18 
  input [18:0] Wgt_1_727, // sfix19_En18 
  input [18:0] Wgt_1_728, // sfix19_En18 
  input [18:0] Wgt_1_729, // sfix19_En18 
  input [18:0] Wgt_1_730, // sfix19_En18 
  input [18:0] Wgt_1_731, // sfix19_En18 
  input [18:0] Wgt_1_732, // sfix19_En18 
  input [18:0] Wgt_1_733, // sfix19_En18 
  input [18:0] Wgt_1_734, // sfix19_En18 
  input [18:0] Wgt_1_735, // sfix19_En18 
  input [18:0] Wgt_1_736, // sfix19_En18 
  input [18:0] Wgt_1_737, // sfix19_En18 
  input [18:0] Wgt_1_738, // sfix19_En18 
  input [18:0] Wgt_1_739, // sfix19_En18 
  input [18:0] Wgt_1_740, // sfix19_En18 
  input [18:0] Wgt_1_741, // sfix19_En18 
  input [18:0] Wgt_1_742, // sfix19_En18 
  input [18:0] Wgt_1_743, // sfix19_En18 
  input [18:0] Wgt_1_744, // sfix19_En18 
  input [18:0] Wgt_1_745, // sfix19_En18 
  input [18:0] Wgt_1_746, // sfix19_En18 
  input [18:0] Wgt_1_747, // sfix19_En18 
  input [18:0] Wgt_1_748, // sfix19_En18 
  input [18:0] Wgt_1_749, // sfix19_En18 
  input [18:0] Wgt_1_750, // sfix19_En18 
  input [18:0] Wgt_1_751, // sfix19_En18 
  input [18:0] Wgt_1_752, // sfix19_En18 
  input [18:0] Wgt_1_753, // sfix19_En18 
  input [18:0] Wgt_1_754, // sfix19_En18 
  input [18:0] Wgt_1_755, // sfix19_En18 
  input [18:0] Wgt_1_756, // sfix19_En18 
  input [18:0] Wgt_1_757, // sfix19_En18 
  input [18:0] Wgt_1_758, // sfix19_En18 
  input [18:0] Wgt_1_759, // sfix19_En18 
  input [18:0] Wgt_1_760, // sfix19_En18 
  input [18:0] Wgt_1_761, // sfix19_En18 
  input [18:0] Wgt_1_762, // sfix19_En18 
  input [18:0] Wgt_1_763, // sfix19_En18 
  input [18:0] Wgt_1_764, // sfix19_En18 
  input [18:0] Wgt_1_765, // sfix19_En18 
  input [18:0] Wgt_1_766, // sfix19_En18 
  input [18:0] Wgt_1_767, // sfix19_En18 
  input [18:0] Wgt_1_768, // sfix19_En18 
  input [18:0] Wgt_1_769, // sfix19_En18 
  input [18:0] Wgt_1_770, // sfix19_En18 
  input [18:0] Wgt_1_771, // sfix19_En18 
  input [18:0] Wgt_1_772, // sfix19_En18 
  input [18:0] Wgt_1_773, // sfix19_En18 
  input [18:0] Wgt_1_774, // sfix19_En18 
  input [18:0] Wgt_1_775, // sfix19_En18 
  input [18:0] Wgt_1_776, // sfix19_En18 
  input [18:0] Wgt_1_777, // sfix19_En18 
  input [18:0] Wgt_1_778, // sfix19_En18 
  input [18:0] Wgt_1_779, // sfix19_En18 
  input [18:0] Wgt_1_780, // sfix19_En18 
  input [18:0] Wgt_1_781, // sfix19_En18 
  input [18:0] Wgt_1_782, // sfix19_En18 
  input [18:0] Wgt_1_783, // sfix19_En18 
  input [18:0] Wgt_1_784, // sfix19_En18 
  input [18:0] Wgt_2_0, // sfix19_En18 
  input [18:0] Wgt_2_1, // sfix19_En18 
  input [18:0] Wgt_2_2, // sfix19_En18 
  input [18:0] Wgt_2_3, // sfix19_En18 
  input [18:0] Wgt_2_4, // sfix19_En18 
  input [18:0] Wgt_2_5, // sfix19_En18 
  input [18:0] Wgt_2_6, // sfix19_En18 
  input [18:0] Wgt_2_7, // sfix19_En18 
  input [18:0] Wgt_2_8, // sfix19_En18 
  input [18:0] Wgt_2_9, // sfix19_En18 
  input [18:0] Wgt_2_10, // sfix19_En18 
  input [18:0] Wgt_2_11, // sfix19_En18 
  input [18:0] Wgt_2_12, // sfix19_En18 
  input [18:0] Wgt_2_13, // sfix19_En18 
  input [18:0] Wgt_2_14, // sfix19_En18 
  input [18:0] Wgt_2_15, // sfix19_En18 
  input [18:0] Wgt_2_16, // sfix19_En18 
  input [18:0] Wgt_2_17, // sfix19_En18 
  input [18:0] Wgt_2_18, // sfix19_En18 
  input [18:0] Wgt_2_19, // sfix19_En18 
  input [18:0] Wgt_2_20, // sfix19_En18 
  input [18:0] Wgt_2_21, // sfix19_En18 
  input [18:0] Wgt_2_22, // sfix19_En18 
  input [18:0] Wgt_2_23, // sfix19_En18 
  input [18:0] Wgt_2_24, // sfix19_En18 
  input [18:0] Wgt_2_25, // sfix19_En18 
  input [18:0] Wgt_2_26, // sfix19_En18 
  input [18:0] Wgt_2_27, // sfix19_En18 
  input [18:0] Wgt_2_28, // sfix19_En18 
  input [18:0] Wgt_2_29, // sfix19_En18 
  input [18:0] Wgt_2_30, // sfix19_En18 
  input [18:0] Wgt_2_31, // sfix19_En18 
  input [18:0] Wgt_2_32, // sfix19_En18 
  input [18:0] Wgt_2_33, // sfix19_En18 
  input [18:0] Wgt_2_34, // sfix19_En18 
  input [18:0] Wgt_2_35, // sfix19_En18 
  input [18:0] Wgt_2_36, // sfix19_En18 
  input [18:0] Wgt_2_37, // sfix19_En18 
  input [18:0] Wgt_2_38, // sfix19_En18 
  input [18:0] Wgt_2_39, // sfix19_En18 
  input [18:0] Wgt_2_40, // sfix19_En18 
  input [18:0] Wgt_2_41, // sfix19_En18 
  input [18:0] Wgt_2_42, // sfix19_En18 
  input [18:0] Wgt_2_43, // sfix19_En18 
  input [18:0] Wgt_2_44, // sfix19_En18 
  input [18:0] Wgt_2_45, // sfix19_En18 
  input [18:0] Wgt_2_46, // sfix19_En18 
  input [18:0] Wgt_2_47, // sfix19_En18 
  input [18:0] Wgt_2_48, // sfix19_En18 
  input [18:0] Wgt_2_49, // sfix19_En18 
  input [18:0] Wgt_2_50, // sfix19_En18 
  input [18:0] Wgt_2_51, // sfix19_En18 
  input [18:0] Wgt_2_52, // sfix19_En18 
  input [18:0] Wgt_2_53, // sfix19_En18 
  input [18:0] Wgt_2_54, // sfix19_En18 
  input [18:0] Wgt_2_55, // sfix19_En18 
  input [18:0] Wgt_2_56, // sfix19_En18 
  input [18:0] Wgt_2_57, // sfix19_En18 
  input [18:0] Wgt_2_58, // sfix19_En18 
  input [18:0] Wgt_2_59, // sfix19_En18 
  input [18:0] Wgt_2_60, // sfix19_En18 
  input [18:0] Wgt_2_61, // sfix19_En18 
  input [18:0] Wgt_2_62, // sfix19_En18 
  input [18:0] Wgt_2_63, // sfix19_En18 
  input [18:0] Wgt_2_64, // sfix19_En18 
  input [18:0] Wgt_2_65, // sfix19_En18 
  input [18:0] Wgt_2_66, // sfix19_En18 
  input [18:0] Wgt_2_67, // sfix19_En18 
  input [18:0] Wgt_2_68, // sfix19_En18 
  input [18:0] Wgt_2_69, // sfix19_En18 
  input [18:0] Wgt_2_70, // sfix19_En18 
  input [18:0] Wgt_2_71, // sfix19_En18 
  input [18:0] Wgt_2_72, // sfix19_En18 
  input [18:0] Wgt_2_73, // sfix19_En18 
  input [18:0] Wgt_2_74, // sfix19_En18 
  input [18:0] Wgt_2_75, // sfix19_En18 
  input [18:0] Wgt_2_76, // sfix19_En18 
  input [18:0] Wgt_2_77, // sfix19_En18 
  input [18:0] Wgt_2_78, // sfix19_En18 
  input [18:0] Wgt_2_79, // sfix19_En18 
  input [18:0] Wgt_2_80, // sfix19_En18 
  input [18:0] Wgt_2_81, // sfix19_En18 
  input [18:0] Wgt_2_82, // sfix19_En18 
  input [18:0] Wgt_2_83, // sfix19_En18 
  input [18:0] Wgt_2_84, // sfix19_En18 
  input [18:0] Wgt_2_85, // sfix19_En18 
  input [18:0] Wgt_2_86, // sfix19_En18 
  input [18:0] Wgt_2_87, // sfix19_En18 
  input [18:0] Wgt_2_88, // sfix19_En18 
  input [18:0] Wgt_2_89, // sfix19_En18 
  input [18:0] Wgt_2_90, // sfix19_En18 
  input [18:0] Wgt_2_91, // sfix19_En18 
  input [18:0] Wgt_2_92, // sfix19_En18 
  input [18:0] Wgt_2_93, // sfix19_En18 
  input [18:0] Wgt_2_94, // sfix19_En18 
  input [18:0] Wgt_2_95, // sfix19_En18 
  input [18:0] Wgt_2_96, // sfix19_En18 
  input [18:0] Wgt_2_97, // sfix19_En18 
  input [18:0] Wgt_2_98, // sfix19_En18 
  input [18:0] Wgt_2_99, // sfix19_En18 
  input [18:0] Wgt_2_100, // sfix19_En18 
  input [18:0] Wgt_2_101, // sfix19_En18 
  input [18:0] Wgt_2_102, // sfix19_En18 
  input [18:0] Wgt_2_103, // sfix19_En18 
  input [18:0] Wgt_2_104, // sfix19_En18 
  input [18:0] Wgt_2_105, // sfix19_En18 
  input [18:0] Wgt_2_106, // sfix19_En18 
  input [18:0] Wgt_2_107, // sfix19_En18 
  input [18:0] Wgt_2_108, // sfix19_En18 
  input [18:0] Wgt_2_109, // sfix19_En18 
  input [18:0] Wgt_2_110, // sfix19_En18 
  input [18:0] Wgt_2_111, // sfix19_En18 
  input [18:0] Wgt_2_112, // sfix19_En18 
  input [18:0] Wgt_2_113, // sfix19_En18 
  input [18:0] Wgt_2_114, // sfix19_En18 
  input [18:0] Wgt_2_115, // sfix19_En18 
  input [18:0] Wgt_2_116, // sfix19_En18 
  input [18:0] Wgt_2_117, // sfix19_En18 
  input [18:0] Wgt_2_118, // sfix19_En18 
  input [18:0] Wgt_2_119, // sfix19_En18 
  input [18:0] Wgt_2_120, // sfix19_En18 
  input [18:0] Wgt_2_121, // sfix19_En18 
  input [18:0] Wgt_2_122, // sfix19_En18 
  input [18:0] Wgt_2_123, // sfix19_En18 
  input [18:0] Wgt_2_124, // sfix19_En18 
  input [18:0] Wgt_2_125, // sfix19_En18 
  input [18:0] Wgt_2_126, // sfix19_En18 
  input [18:0] Wgt_2_127, // sfix19_En18 
  input [18:0] Wgt_2_128, // sfix19_En18 
  input [18:0] Wgt_2_129, // sfix19_En18 
  input [18:0] Wgt_2_130, // sfix19_En18 
  input [18:0] Wgt_2_131, // sfix19_En18 
  input [18:0] Wgt_2_132, // sfix19_En18 
  input [18:0] Wgt_2_133, // sfix19_En18 
  input [18:0] Wgt_2_134, // sfix19_En18 
  input [18:0] Wgt_2_135, // sfix19_En18 
  input [18:0] Wgt_2_136, // sfix19_En18 
  input [18:0] Wgt_2_137, // sfix19_En18 
  input [18:0] Wgt_2_138, // sfix19_En18 
  input [18:0] Wgt_2_139, // sfix19_En18 
  input [18:0] Wgt_2_140, // sfix19_En18 
  input [18:0] Wgt_2_141, // sfix19_En18 
  input [18:0] Wgt_2_142, // sfix19_En18 
  input [18:0] Wgt_2_143, // sfix19_En18 
  input [18:0] Wgt_2_144, // sfix19_En18 
  input [18:0] Wgt_2_145, // sfix19_En18 
  input [18:0] Wgt_2_146, // sfix19_En18 
  input [18:0] Wgt_2_147, // sfix19_En18 
  input [18:0] Wgt_2_148, // sfix19_En18 
  input [18:0] Wgt_2_149, // sfix19_En18 
  input [18:0] Wgt_2_150, // sfix19_En18 
  input [18:0] Wgt_2_151, // sfix19_En18 
  input [18:0] Wgt_2_152, // sfix19_En18 
  input [18:0] Wgt_2_153, // sfix19_En18 
  input [18:0] Wgt_2_154, // sfix19_En18 
  input [18:0] Wgt_2_155, // sfix19_En18 
  input [18:0] Wgt_2_156, // sfix19_En18 
  input [18:0] Wgt_2_157, // sfix19_En18 
  input [18:0] Wgt_2_158, // sfix19_En18 
  input [18:0] Wgt_2_159, // sfix19_En18 
  input [18:0] Wgt_2_160, // sfix19_En18 
  input [18:0] Wgt_2_161, // sfix19_En18 
  input [18:0] Wgt_2_162, // sfix19_En18 
  input [18:0] Wgt_2_163, // sfix19_En18 
  input [18:0] Wgt_2_164, // sfix19_En18 
  input [18:0] Wgt_2_165, // sfix19_En18 
  input [18:0] Wgt_2_166, // sfix19_En18 
  input [18:0] Wgt_2_167, // sfix19_En18 
  input [18:0] Wgt_2_168, // sfix19_En18 
  input [18:0] Wgt_2_169, // sfix19_En18 
  input [18:0] Wgt_2_170, // sfix19_En18 
  input [18:0] Wgt_2_171, // sfix19_En18 
  input [18:0] Wgt_2_172, // sfix19_En18 
  input [18:0] Wgt_2_173, // sfix19_En18 
  input [18:0] Wgt_2_174, // sfix19_En18 
  input [18:0] Wgt_2_175, // sfix19_En18 
  input [18:0] Wgt_2_176, // sfix19_En18 
  input [18:0] Wgt_2_177, // sfix19_En18 
  input [18:0] Wgt_2_178, // sfix19_En18 
  input [18:0] Wgt_2_179, // sfix19_En18 
  input [18:0] Wgt_2_180, // sfix19_En18 
  input [18:0] Wgt_2_181, // sfix19_En18 
  input [18:0] Wgt_2_182, // sfix19_En18 
  input [18:0] Wgt_2_183, // sfix19_En18 
  input [18:0] Wgt_2_184, // sfix19_En18 
  input [18:0] Wgt_2_185, // sfix19_En18 
  input [18:0] Wgt_2_186, // sfix19_En18 
  input [18:0] Wgt_2_187, // sfix19_En18 
  input [18:0] Wgt_2_188, // sfix19_En18 
  input [18:0] Wgt_2_189, // sfix19_En18 
  input [18:0] Wgt_2_190, // sfix19_En18 
  input [18:0] Wgt_2_191, // sfix19_En18 
  input [18:0] Wgt_2_192, // sfix19_En18 
  input [18:0] Wgt_2_193, // sfix19_En18 
  input [18:0] Wgt_2_194, // sfix19_En18 
  input [18:0] Wgt_2_195, // sfix19_En18 
  input [18:0] Wgt_2_196, // sfix19_En18 
  input [18:0] Wgt_2_197, // sfix19_En18 
  input [18:0] Wgt_2_198, // sfix19_En18 
  input [18:0] Wgt_2_199, // sfix19_En18 
  input [18:0] Wgt_2_200, // sfix19_En18 
  input [18:0] Wgt_2_201, // sfix19_En18 
  input [18:0] Wgt_2_202, // sfix19_En18 
  input [18:0] Wgt_2_203, // sfix19_En18 
  input [18:0] Wgt_2_204, // sfix19_En18 
  input [18:0] Wgt_2_205, // sfix19_En18 
  input [18:0] Wgt_2_206, // sfix19_En18 
  input [18:0] Wgt_2_207, // sfix19_En18 
  input [18:0] Wgt_2_208, // sfix19_En18 
  input [18:0] Wgt_2_209, // sfix19_En18 
  input [18:0] Wgt_2_210, // sfix19_En18 
  input [18:0] Wgt_2_211, // sfix19_En18 
  input [18:0] Wgt_2_212, // sfix19_En18 
  input [18:0] Wgt_2_213, // sfix19_En18 
  input [18:0] Wgt_2_214, // sfix19_En18 
  input [18:0] Wgt_2_215, // sfix19_En18 
  input [18:0] Wgt_2_216, // sfix19_En18 
  input [18:0] Wgt_2_217, // sfix19_En18 
  input [18:0] Wgt_2_218, // sfix19_En18 
  input [18:0] Wgt_2_219, // sfix19_En18 
  input [18:0] Wgt_2_220, // sfix19_En18 
  input [18:0] Wgt_2_221, // sfix19_En18 
  input [18:0] Wgt_2_222, // sfix19_En18 
  input [18:0] Wgt_2_223, // sfix19_En18 
  input [18:0] Wgt_2_224, // sfix19_En18 
  input [18:0] Wgt_2_225, // sfix19_En18 
  input [18:0] Wgt_2_226, // sfix19_En18 
  input [18:0] Wgt_2_227, // sfix19_En18 
  input [18:0] Wgt_2_228, // sfix19_En18 
  input [18:0] Wgt_2_229, // sfix19_En18 
  input [18:0] Wgt_2_230, // sfix19_En18 
  input [18:0] Wgt_2_231, // sfix19_En18 
  input [18:0] Wgt_2_232, // sfix19_En18 
  input [18:0] Wgt_2_233, // sfix19_En18 
  input [18:0] Wgt_2_234, // sfix19_En18 
  input [18:0] Wgt_2_235, // sfix19_En18 
  input [18:0] Wgt_2_236, // sfix19_En18 
  input [18:0] Wgt_2_237, // sfix19_En18 
  input [18:0] Wgt_2_238, // sfix19_En18 
  input [18:0] Wgt_2_239, // sfix19_En18 
  input [18:0] Wgt_2_240, // sfix19_En18 
  input [18:0] Wgt_2_241, // sfix19_En18 
  input [18:0] Wgt_2_242, // sfix19_En18 
  input [18:0] Wgt_2_243, // sfix19_En18 
  input [18:0] Wgt_2_244, // sfix19_En18 
  input [18:0] Wgt_2_245, // sfix19_En18 
  input [18:0] Wgt_2_246, // sfix19_En18 
  input [18:0] Wgt_2_247, // sfix19_En18 
  input [18:0] Wgt_2_248, // sfix19_En18 
  input [18:0] Wgt_2_249, // sfix19_En18 
  input [18:0] Wgt_2_250, // sfix19_En18 
  input [18:0] Wgt_2_251, // sfix19_En18 
  input [18:0] Wgt_2_252, // sfix19_En18 
  input [18:0] Wgt_2_253, // sfix19_En18 
  input [18:0] Wgt_2_254, // sfix19_En18 
  input [18:0] Wgt_2_255, // sfix19_En18 
  input [18:0] Wgt_2_256, // sfix19_En18 
  input [18:0] Wgt_2_257, // sfix19_En18 
  input [18:0] Wgt_2_258, // sfix19_En18 
  input [18:0] Wgt_2_259, // sfix19_En18 
  input [18:0] Wgt_2_260, // sfix19_En18 
  input [18:0] Wgt_2_261, // sfix19_En18 
  input [18:0] Wgt_2_262, // sfix19_En18 
  input [18:0] Wgt_2_263, // sfix19_En18 
  input [18:0] Wgt_2_264, // sfix19_En18 
  input [18:0] Wgt_2_265, // sfix19_En18 
  input [18:0] Wgt_2_266, // sfix19_En18 
  input [18:0] Wgt_2_267, // sfix19_En18 
  input [18:0] Wgt_2_268, // sfix19_En18 
  input [18:0] Wgt_2_269, // sfix19_En18 
  input [18:0] Wgt_2_270, // sfix19_En18 
  input [18:0] Wgt_2_271, // sfix19_En18 
  input [18:0] Wgt_2_272, // sfix19_En18 
  input [18:0] Wgt_2_273, // sfix19_En18 
  input [18:0] Wgt_2_274, // sfix19_En18 
  input [18:0] Wgt_2_275, // sfix19_En18 
  input [18:0] Wgt_2_276, // sfix19_En18 
  input [18:0] Wgt_2_277, // sfix19_En18 
  input [18:0] Wgt_2_278, // sfix19_En18 
  input [18:0] Wgt_2_279, // sfix19_En18 
  input [18:0] Wgt_2_280, // sfix19_En18 
  input [18:0] Wgt_2_281, // sfix19_En18 
  input [18:0] Wgt_2_282, // sfix19_En18 
  input [18:0] Wgt_2_283, // sfix19_En18 
  input [18:0] Wgt_2_284, // sfix19_En18 
  input [18:0] Wgt_2_285, // sfix19_En18 
  input [18:0] Wgt_2_286, // sfix19_En18 
  input [18:0] Wgt_2_287, // sfix19_En18 
  input [18:0] Wgt_2_288, // sfix19_En18 
  input [18:0] Wgt_2_289, // sfix19_En18 
  input [18:0] Wgt_2_290, // sfix19_En18 
  input [18:0] Wgt_2_291, // sfix19_En18 
  input [18:0] Wgt_2_292, // sfix19_En18 
  input [18:0] Wgt_2_293, // sfix19_En18 
  input [18:0] Wgt_2_294, // sfix19_En18 
  input [18:0] Wgt_2_295, // sfix19_En18 
  input [18:0] Wgt_2_296, // sfix19_En18 
  input [18:0] Wgt_2_297, // sfix19_En18 
  input [18:0] Wgt_2_298, // sfix19_En18 
  input [18:0] Wgt_2_299, // sfix19_En18 
  input [18:0] Wgt_2_300, // sfix19_En18 
  input [18:0] Wgt_2_301, // sfix19_En18 
  input [18:0] Wgt_2_302, // sfix19_En18 
  input [18:0] Wgt_2_303, // sfix19_En18 
  input [18:0] Wgt_2_304, // sfix19_En18 
  input [18:0] Wgt_2_305, // sfix19_En18 
  input [18:0] Wgt_2_306, // sfix19_En18 
  input [18:0] Wgt_2_307, // sfix19_En18 
  input [18:0] Wgt_2_308, // sfix19_En18 
  input [18:0] Wgt_2_309, // sfix19_En18 
  input [18:0] Wgt_2_310, // sfix19_En18 
  input [18:0] Wgt_2_311, // sfix19_En18 
  input [18:0] Wgt_2_312, // sfix19_En18 
  input [18:0] Wgt_2_313, // sfix19_En18 
  input [18:0] Wgt_2_314, // sfix19_En18 
  input [18:0] Wgt_2_315, // sfix19_En18 
  input [18:0] Wgt_2_316, // sfix19_En18 
  input [18:0] Wgt_2_317, // sfix19_En18 
  input [18:0] Wgt_2_318, // sfix19_En18 
  input [18:0] Wgt_2_319, // sfix19_En18 
  input [18:0] Wgt_2_320, // sfix19_En18 
  input [18:0] Wgt_2_321, // sfix19_En18 
  input [18:0] Wgt_2_322, // sfix19_En18 
  input [18:0] Wgt_2_323, // sfix19_En18 
  input [18:0] Wgt_2_324, // sfix19_En18 
  input [18:0] Wgt_2_325, // sfix19_En18 
  input [18:0] Wgt_2_326, // sfix19_En18 
  input [18:0] Wgt_2_327, // sfix19_En18 
  input [18:0] Wgt_2_328, // sfix19_En18 
  input [18:0] Wgt_2_329, // sfix19_En18 
  input [18:0] Wgt_2_330, // sfix19_En18 
  input [18:0] Wgt_2_331, // sfix19_En18 
  input [18:0] Wgt_2_332, // sfix19_En18 
  input [18:0] Wgt_2_333, // sfix19_En18 
  input [18:0] Wgt_2_334, // sfix19_En18 
  input [18:0] Wgt_2_335, // sfix19_En18 
  input [18:0] Wgt_2_336, // sfix19_En18 
  input [18:0] Wgt_2_337, // sfix19_En18 
  input [18:0] Wgt_2_338, // sfix19_En18 
  input [18:0] Wgt_2_339, // sfix19_En18 
  input [18:0] Wgt_2_340, // sfix19_En18 
  input [18:0] Wgt_2_341, // sfix19_En18 
  input [18:0] Wgt_2_342, // sfix19_En18 
  input [18:0] Wgt_2_343, // sfix19_En18 
  input [18:0] Wgt_2_344, // sfix19_En18 
  input [18:0] Wgt_2_345, // sfix19_En18 
  input [18:0] Wgt_2_346, // sfix19_En18 
  input [18:0] Wgt_2_347, // sfix19_En18 
  input [18:0] Wgt_2_348, // sfix19_En18 
  input [18:0] Wgt_2_349, // sfix19_En18 
  input [18:0] Wgt_2_350, // sfix19_En18 
  input [18:0] Wgt_2_351, // sfix19_En18 
  input [18:0] Wgt_2_352, // sfix19_En18 
  input [18:0] Wgt_2_353, // sfix19_En18 
  input [18:0] Wgt_2_354, // sfix19_En18 
  input [18:0] Wgt_2_355, // sfix19_En18 
  input [18:0] Wgt_2_356, // sfix19_En18 
  input [18:0] Wgt_2_357, // sfix19_En18 
  input [18:0] Wgt_2_358, // sfix19_En18 
  input [18:0] Wgt_2_359, // sfix19_En18 
  input [18:0] Wgt_2_360, // sfix19_En18 
  input [18:0] Wgt_2_361, // sfix19_En18 
  input [18:0] Wgt_2_362, // sfix19_En18 
  input [18:0] Wgt_2_363, // sfix19_En18 
  input [18:0] Wgt_2_364, // sfix19_En18 
  input [18:0] Wgt_2_365, // sfix19_En18 
  input [18:0] Wgt_2_366, // sfix19_En18 
  input [18:0] Wgt_2_367, // sfix19_En18 
  input [18:0] Wgt_2_368, // sfix19_En18 
  input [18:0] Wgt_2_369, // sfix19_En18 
  input [18:0] Wgt_2_370, // sfix19_En18 
  input [18:0] Wgt_2_371, // sfix19_En18 
  input [18:0] Wgt_2_372, // sfix19_En18 
  input [18:0] Wgt_2_373, // sfix19_En18 
  input [18:0] Wgt_2_374, // sfix19_En18 
  input [18:0] Wgt_2_375, // sfix19_En18 
  input [18:0] Wgt_2_376, // sfix19_En18 
  input [18:0] Wgt_2_377, // sfix19_En18 
  input [18:0] Wgt_2_378, // sfix19_En18 
  input [18:0] Wgt_2_379, // sfix19_En18 
  input [18:0] Wgt_2_380, // sfix19_En18 
  input [18:0] Wgt_2_381, // sfix19_En18 
  input [18:0] Wgt_2_382, // sfix19_En18 
  input [18:0] Wgt_2_383, // sfix19_En18 
  input [18:0] Wgt_2_384, // sfix19_En18 
  input [18:0] Wgt_2_385, // sfix19_En18 
  input [18:0] Wgt_2_386, // sfix19_En18 
  input [18:0] Wgt_2_387, // sfix19_En18 
  input [18:0] Wgt_2_388, // sfix19_En18 
  input [18:0] Wgt_2_389, // sfix19_En18 
  input [18:0] Wgt_2_390, // sfix19_En18 
  input [18:0] Wgt_2_391, // sfix19_En18 
  input [18:0] Wgt_2_392, // sfix19_En18 
  input [18:0] Wgt_2_393, // sfix19_En18 
  input [18:0] Wgt_2_394, // sfix19_En18 
  input [18:0] Wgt_2_395, // sfix19_En18 
  input [18:0] Wgt_2_396, // sfix19_En18 
  input [18:0] Wgt_2_397, // sfix19_En18 
  input [18:0] Wgt_2_398, // sfix19_En18 
  input [18:0] Wgt_2_399, // sfix19_En18 
  input [18:0] Wgt_2_400, // sfix19_En18 
  input [18:0] Wgt_2_401, // sfix19_En18 
  input [18:0] Wgt_2_402, // sfix19_En18 
  input [18:0] Wgt_2_403, // sfix19_En18 
  input [18:0] Wgt_2_404, // sfix19_En18 
  input [18:0] Wgt_2_405, // sfix19_En18 
  input [18:0] Wgt_2_406, // sfix19_En18 
  input [18:0] Wgt_2_407, // sfix19_En18 
  input [18:0] Wgt_2_408, // sfix19_En18 
  input [18:0] Wgt_2_409, // sfix19_En18 
  input [18:0] Wgt_2_410, // sfix19_En18 
  input [18:0] Wgt_2_411, // sfix19_En18 
  input [18:0] Wgt_2_412, // sfix19_En18 
  input [18:0] Wgt_2_413, // sfix19_En18 
  input [18:0] Wgt_2_414, // sfix19_En18 
  input [18:0] Wgt_2_415, // sfix19_En18 
  input [18:0] Wgt_2_416, // sfix19_En18 
  input [18:0] Wgt_2_417, // sfix19_En18 
  input [18:0] Wgt_2_418, // sfix19_En18 
  input [18:0] Wgt_2_419, // sfix19_En18 
  input [18:0] Wgt_2_420, // sfix19_En18 
  input [18:0] Wgt_2_421, // sfix19_En18 
  input [18:0] Wgt_2_422, // sfix19_En18 
  input [18:0] Wgt_2_423, // sfix19_En18 
  input [18:0] Wgt_2_424, // sfix19_En18 
  input [18:0] Wgt_2_425, // sfix19_En18 
  input [18:0] Wgt_2_426, // sfix19_En18 
  input [18:0] Wgt_2_427, // sfix19_En18 
  input [18:0] Wgt_2_428, // sfix19_En18 
  input [18:0] Wgt_2_429, // sfix19_En18 
  input [18:0] Wgt_2_430, // sfix19_En18 
  input [18:0] Wgt_2_431, // sfix19_En18 
  input [18:0] Wgt_2_432, // sfix19_En18 
  input [18:0] Wgt_2_433, // sfix19_En18 
  input [18:0] Wgt_2_434, // sfix19_En18 
  input [18:0] Wgt_2_435, // sfix19_En18 
  input [18:0] Wgt_2_436, // sfix19_En18 
  input [18:0] Wgt_2_437, // sfix19_En18 
  input [18:0] Wgt_2_438, // sfix19_En18 
  input [18:0] Wgt_2_439, // sfix19_En18 
  input [18:0] Wgt_2_440, // sfix19_En18 
  input [18:0] Wgt_2_441, // sfix19_En18 
  input [18:0] Wgt_2_442, // sfix19_En18 
  input [18:0] Wgt_2_443, // sfix19_En18 
  input [18:0] Wgt_2_444, // sfix19_En18 
  input [18:0] Wgt_2_445, // sfix19_En18 
  input [18:0] Wgt_2_446, // sfix19_En18 
  input [18:0] Wgt_2_447, // sfix19_En18 
  input [18:0] Wgt_2_448, // sfix19_En18 
  input [18:0] Wgt_2_449, // sfix19_En18 
  input [18:0] Wgt_2_450, // sfix19_En18 
  input [18:0] Wgt_2_451, // sfix19_En18 
  input [18:0] Wgt_2_452, // sfix19_En18 
  input [18:0] Wgt_2_453, // sfix19_En18 
  input [18:0] Wgt_2_454, // sfix19_En18 
  input [18:0] Wgt_2_455, // sfix19_En18 
  input [18:0] Wgt_2_456, // sfix19_En18 
  input [18:0] Wgt_2_457, // sfix19_En18 
  input [18:0] Wgt_2_458, // sfix19_En18 
  input [18:0] Wgt_2_459, // sfix19_En18 
  input [18:0] Wgt_2_460, // sfix19_En18 
  input [18:0] Wgt_2_461, // sfix19_En18 
  input [18:0] Wgt_2_462, // sfix19_En18 
  input [18:0] Wgt_2_463, // sfix19_En18 
  input [18:0] Wgt_2_464, // sfix19_En18 
  input [18:0] Wgt_2_465, // sfix19_En18 
  input [18:0] Wgt_2_466, // sfix19_En18 
  input [18:0] Wgt_2_467, // sfix19_En18 
  input [18:0] Wgt_2_468, // sfix19_En18 
  input [18:0] Wgt_2_469, // sfix19_En18 
  input [18:0] Wgt_2_470, // sfix19_En18 
  input [18:0] Wgt_2_471, // sfix19_En18 
  input [18:0] Wgt_2_472, // sfix19_En18 
  input [18:0] Wgt_2_473, // sfix19_En18 
  input [18:0] Wgt_2_474, // sfix19_En18 
  input [18:0] Wgt_2_475, // sfix19_En18 
  input [18:0] Wgt_2_476, // sfix19_En18 
  input [18:0] Wgt_2_477, // sfix19_En18 
  input [18:0] Wgt_2_478, // sfix19_En18 
  input [18:0] Wgt_2_479, // sfix19_En18 
  input [18:0] Wgt_2_480, // sfix19_En18 
  input [18:0] Wgt_2_481, // sfix19_En18 
  input [18:0] Wgt_2_482, // sfix19_En18 
  input [18:0] Wgt_2_483, // sfix19_En18 
  input [18:0] Wgt_2_484, // sfix19_En18 
  input [18:0] Wgt_2_485, // sfix19_En18 
  input [18:0] Wgt_2_486, // sfix19_En18 
  input [18:0] Wgt_2_487, // sfix19_En18 
  input [18:0] Wgt_2_488, // sfix19_En18 
  input [18:0] Wgt_2_489, // sfix19_En18 
  input [18:0] Wgt_2_490, // sfix19_En18 
  input [18:0] Wgt_2_491, // sfix19_En18 
  input [18:0] Wgt_2_492, // sfix19_En18 
  input [18:0] Wgt_2_493, // sfix19_En18 
  input [18:0] Wgt_2_494, // sfix19_En18 
  input [18:0] Wgt_2_495, // sfix19_En18 
  input [18:0] Wgt_2_496, // sfix19_En18 
  input [18:0] Wgt_2_497, // sfix19_En18 
  input [18:0] Wgt_2_498, // sfix19_En18 
  input [18:0] Wgt_2_499, // sfix19_En18 
  input [18:0] Wgt_2_500, // sfix19_En18 
  input [18:0] Wgt_2_501, // sfix19_En18 
  input [18:0] Wgt_2_502, // sfix19_En18 
  input [18:0] Wgt_2_503, // sfix19_En18 
  input [18:0] Wgt_2_504, // sfix19_En18 
  input [18:0] Wgt_2_505, // sfix19_En18 
  input [18:0] Wgt_2_506, // sfix19_En18 
  input [18:0] Wgt_2_507, // sfix19_En18 
  input [18:0] Wgt_2_508, // sfix19_En18 
  input [18:0] Wgt_2_509, // sfix19_En18 
  input [18:0] Wgt_2_510, // sfix19_En18 
  input [18:0] Wgt_2_511, // sfix19_En18 
  input [18:0] Wgt_2_512, // sfix19_En18 
  input [18:0] Wgt_2_513, // sfix19_En18 
  input [18:0] Wgt_2_514, // sfix19_En18 
  input [18:0] Wgt_2_515, // sfix19_En18 
  input [18:0] Wgt_2_516, // sfix19_En18 
  input [18:0] Wgt_2_517, // sfix19_En18 
  input [18:0] Wgt_2_518, // sfix19_En18 
  input [18:0] Wgt_2_519, // sfix19_En18 
  input [18:0] Wgt_2_520, // sfix19_En18 
  input [18:0] Wgt_2_521, // sfix19_En18 
  input [18:0] Wgt_2_522, // sfix19_En18 
  input [18:0] Wgt_2_523, // sfix19_En18 
  input [18:0] Wgt_2_524, // sfix19_En18 
  input [18:0] Wgt_2_525, // sfix19_En18 
  input [18:0] Wgt_2_526, // sfix19_En18 
  input [18:0] Wgt_2_527, // sfix19_En18 
  input [18:0] Wgt_2_528, // sfix19_En18 
  input [18:0] Wgt_2_529, // sfix19_En18 
  input [18:0] Wgt_2_530, // sfix19_En18 
  input [18:0] Wgt_2_531, // sfix19_En18 
  input [18:0] Wgt_2_532, // sfix19_En18 
  input [18:0] Wgt_2_533, // sfix19_En18 
  input [18:0] Wgt_2_534, // sfix19_En18 
  input [18:0] Wgt_2_535, // sfix19_En18 
  input [18:0] Wgt_2_536, // sfix19_En18 
  input [18:0] Wgt_2_537, // sfix19_En18 
  input [18:0] Wgt_2_538, // sfix19_En18 
  input [18:0] Wgt_2_539, // sfix19_En18 
  input [18:0] Wgt_2_540, // sfix19_En18 
  input [18:0] Wgt_2_541, // sfix19_En18 
  input [18:0] Wgt_2_542, // sfix19_En18 
  input [18:0] Wgt_2_543, // sfix19_En18 
  input [18:0] Wgt_2_544, // sfix19_En18 
  input [18:0] Wgt_2_545, // sfix19_En18 
  input [18:0] Wgt_2_546, // sfix19_En18 
  input [18:0] Wgt_2_547, // sfix19_En18 
  input [18:0] Wgt_2_548, // sfix19_En18 
  input [18:0] Wgt_2_549, // sfix19_En18 
  input [18:0] Wgt_2_550, // sfix19_En18 
  input [18:0] Wgt_2_551, // sfix19_En18 
  input [18:0] Wgt_2_552, // sfix19_En18 
  input [18:0] Wgt_2_553, // sfix19_En18 
  input [18:0] Wgt_2_554, // sfix19_En18 
  input [18:0] Wgt_2_555, // sfix19_En18 
  input [18:0] Wgt_2_556, // sfix19_En18 
  input [18:0] Wgt_2_557, // sfix19_En18 
  input [18:0] Wgt_2_558, // sfix19_En18 
  input [18:0] Wgt_2_559, // sfix19_En18 
  input [18:0] Wgt_2_560, // sfix19_En18 
  input [18:0] Wgt_2_561, // sfix19_En18 
  input [18:0] Wgt_2_562, // sfix19_En18 
  input [18:0] Wgt_2_563, // sfix19_En18 
  input [18:0] Wgt_2_564, // sfix19_En18 
  input [18:0] Wgt_2_565, // sfix19_En18 
  input [18:0] Wgt_2_566, // sfix19_En18 
  input [18:0] Wgt_2_567, // sfix19_En18 
  input [18:0] Wgt_2_568, // sfix19_En18 
  input [18:0] Wgt_2_569, // sfix19_En18 
  input [18:0] Wgt_2_570, // sfix19_En18 
  input [18:0] Wgt_2_571, // sfix19_En18 
  input [18:0] Wgt_2_572, // sfix19_En18 
  input [18:0] Wgt_2_573, // sfix19_En18 
  input [18:0] Wgt_2_574, // sfix19_En18 
  input [18:0] Wgt_2_575, // sfix19_En18 
  input [18:0] Wgt_2_576, // sfix19_En18 
  input [18:0] Wgt_2_577, // sfix19_En18 
  input [18:0] Wgt_2_578, // sfix19_En18 
  input [18:0] Wgt_2_579, // sfix19_En18 
  input [18:0] Wgt_2_580, // sfix19_En18 
  input [18:0] Wgt_2_581, // sfix19_En18 
  input [18:0] Wgt_2_582, // sfix19_En18 
  input [18:0] Wgt_2_583, // sfix19_En18 
  input [18:0] Wgt_2_584, // sfix19_En18 
  input [18:0] Wgt_2_585, // sfix19_En18 
  input [18:0] Wgt_2_586, // sfix19_En18 
  input [18:0] Wgt_2_587, // sfix19_En18 
  input [18:0] Wgt_2_588, // sfix19_En18 
  input [18:0] Wgt_2_589, // sfix19_En18 
  input [18:0] Wgt_2_590, // sfix19_En18 
  input [18:0] Wgt_2_591, // sfix19_En18 
  input [18:0] Wgt_2_592, // sfix19_En18 
  input [18:0] Wgt_2_593, // sfix19_En18 
  input [18:0] Wgt_2_594, // sfix19_En18 
  input [18:0] Wgt_2_595, // sfix19_En18 
  input [18:0] Wgt_2_596, // sfix19_En18 
  input [18:0] Wgt_2_597, // sfix19_En18 
  input [18:0] Wgt_2_598, // sfix19_En18 
  input [18:0] Wgt_2_599, // sfix19_En18 
  input [18:0] Wgt_2_600, // sfix19_En18 
  input [18:0] Wgt_2_601, // sfix19_En18 
  input [18:0] Wgt_2_602, // sfix19_En18 
  input [18:0] Wgt_2_603, // sfix19_En18 
  input [18:0] Wgt_2_604, // sfix19_En18 
  input [18:0] Wgt_2_605, // sfix19_En18 
  input [18:0] Wgt_2_606, // sfix19_En18 
  input [18:0] Wgt_2_607, // sfix19_En18 
  input [18:0] Wgt_2_608, // sfix19_En18 
  input [18:0] Wgt_2_609, // sfix19_En18 
  input [18:0] Wgt_2_610, // sfix19_En18 
  input [18:0] Wgt_2_611, // sfix19_En18 
  input [18:0] Wgt_2_612, // sfix19_En18 
  input [18:0] Wgt_2_613, // sfix19_En18 
  input [18:0] Wgt_2_614, // sfix19_En18 
  input [18:0] Wgt_2_615, // sfix19_En18 
  input [18:0] Wgt_2_616, // sfix19_En18 
  input [18:0] Wgt_2_617, // sfix19_En18 
  input [18:0] Wgt_2_618, // sfix19_En18 
  input [18:0] Wgt_2_619, // sfix19_En18 
  input [18:0] Wgt_2_620, // sfix19_En18 
  input [18:0] Wgt_2_621, // sfix19_En18 
  input [18:0] Wgt_2_622, // sfix19_En18 
  input [18:0] Wgt_2_623, // sfix19_En18 
  input [18:0] Wgt_2_624, // sfix19_En18 
  input [18:0] Wgt_2_625, // sfix19_En18 
  input [18:0] Wgt_2_626, // sfix19_En18 
  input [18:0] Wgt_2_627, // sfix19_En18 
  input [18:0] Wgt_2_628, // sfix19_En18 
  input [18:0] Wgt_2_629, // sfix19_En18 
  input [18:0] Wgt_2_630, // sfix19_En18 
  input [18:0] Wgt_2_631, // sfix19_En18 
  input [18:0] Wgt_2_632, // sfix19_En18 
  input [18:0] Wgt_2_633, // sfix19_En18 
  input [18:0] Wgt_2_634, // sfix19_En18 
  input [18:0] Wgt_2_635, // sfix19_En18 
  input [18:0] Wgt_2_636, // sfix19_En18 
  input [18:0] Wgt_2_637, // sfix19_En18 
  input [18:0] Wgt_2_638, // sfix19_En18 
  input [18:0] Wgt_2_639, // sfix19_En18 
  input [18:0] Wgt_2_640, // sfix19_En18 
  input [18:0] Wgt_2_641, // sfix19_En18 
  input [18:0] Wgt_2_642, // sfix19_En18 
  input [18:0] Wgt_2_643, // sfix19_En18 
  input [18:0] Wgt_2_644, // sfix19_En18 
  input [18:0] Wgt_2_645, // sfix19_En18 
  input [18:0] Wgt_2_646, // sfix19_En18 
  input [18:0] Wgt_2_647, // sfix19_En18 
  input [18:0] Wgt_2_648, // sfix19_En18 
  input [18:0] Wgt_2_649, // sfix19_En18 
  input [18:0] Wgt_2_650, // sfix19_En18 
  input [18:0] Wgt_2_651, // sfix19_En18 
  input [18:0] Wgt_2_652, // sfix19_En18 
  input [18:0] Wgt_2_653, // sfix19_En18 
  input [18:0] Wgt_2_654, // sfix19_En18 
  input [18:0] Wgt_2_655, // sfix19_En18 
  input [18:0] Wgt_2_656, // sfix19_En18 
  input [18:0] Wgt_2_657, // sfix19_En18 
  input [18:0] Wgt_2_658, // sfix19_En18 
  input [18:0] Wgt_2_659, // sfix19_En18 
  input [18:0] Wgt_2_660, // sfix19_En18 
  input [18:0] Wgt_2_661, // sfix19_En18 
  input [18:0] Wgt_2_662, // sfix19_En18 
  input [18:0] Wgt_2_663, // sfix19_En18 
  input [18:0] Wgt_2_664, // sfix19_En18 
  input [18:0] Wgt_2_665, // sfix19_En18 
  input [18:0] Wgt_2_666, // sfix19_En18 
  input [18:0] Wgt_2_667, // sfix19_En18 
  input [18:0] Wgt_2_668, // sfix19_En18 
  input [18:0] Wgt_2_669, // sfix19_En18 
  input [18:0] Wgt_2_670, // sfix19_En18 
  input [18:0] Wgt_2_671, // sfix19_En18 
  input [18:0] Wgt_2_672, // sfix19_En18 
  input [18:0] Wgt_2_673, // sfix19_En18 
  input [18:0] Wgt_2_674, // sfix19_En18 
  input [18:0] Wgt_2_675, // sfix19_En18 
  input [18:0] Wgt_2_676, // sfix19_En18 
  input [18:0] Wgt_2_677, // sfix19_En18 
  input [18:0] Wgt_2_678, // sfix19_En18 
  input [18:0] Wgt_2_679, // sfix19_En18 
  input [18:0] Wgt_2_680, // sfix19_En18 
  input [18:0] Wgt_2_681, // sfix19_En18 
  input [18:0] Wgt_2_682, // sfix19_En18 
  input [18:0] Wgt_2_683, // sfix19_En18 
  input [18:0] Wgt_2_684, // sfix19_En18 
  input [18:0] Wgt_2_685, // sfix19_En18 
  input [18:0] Wgt_2_686, // sfix19_En18 
  input [18:0] Wgt_2_687, // sfix19_En18 
  input [18:0] Wgt_2_688, // sfix19_En18 
  input [18:0] Wgt_2_689, // sfix19_En18 
  input [18:0] Wgt_2_690, // sfix19_En18 
  input [18:0] Wgt_2_691, // sfix19_En18 
  input [18:0] Wgt_2_692, // sfix19_En18 
  input [18:0] Wgt_2_693, // sfix19_En18 
  input [18:0] Wgt_2_694, // sfix19_En18 
  input [18:0] Wgt_2_695, // sfix19_En18 
  input [18:0] Wgt_2_696, // sfix19_En18 
  input [18:0] Wgt_2_697, // sfix19_En18 
  input [18:0] Wgt_2_698, // sfix19_En18 
  input [18:0] Wgt_2_699, // sfix19_En18 
  input [18:0] Wgt_2_700, // sfix19_En18 
  input [18:0] Wgt_2_701, // sfix19_En18 
  input [18:0] Wgt_2_702, // sfix19_En18 
  input [18:0] Wgt_2_703, // sfix19_En18 
  input [18:0] Wgt_2_704, // sfix19_En18 
  input [18:0] Wgt_2_705, // sfix19_En18 
  input [18:0] Wgt_2_706, // sfix19_En18 
  input [18:0] Wgt_2_707, // sfix19_En18 
  input [18:0] Wgt_2_708, // sfix19_En18 
  input [18:0] Wgt_2_709, // sfix19_En18 
  input [18:0] Wgt_2_710, // sfix19_En18 
  input [18:0] Wgt_2_711, // sfix19_En18 
  input [18:0] Wgt_2_712, // sfix19_En18 
  input [18:0] Wgt_2_713, // sfix19_En18 
  input [18:0] Wgt_2_714, // sfix19_En18 
  input [18:0] Wgt_2_715, // sfix19_En18 
  input [18:0] Wgt_2_716, // sfix19_En18 
  input [18:0] Wgt_2_717, // sfix19_En18 
  input [18:0] Wgt_2_718, // sfix19_En18 
  input [18:0] Wgt_2_719, // sfix19_En18 
  input [18:0] Wgt_2_720, // sfix19_En18 
  input [18:0] Wgt_2_721, // sfix19_En18 
  input [18:0] Wgt_2_722, // sfix19_En18 
  input [18:0] Wgt_2_723, // sfix19_En18 
  input [18:0] Wgt_2_724, // sfix19_En18 
  input [18:0] Wgt_2_725, // sfix19_En18 
  input [18:0] Wgt_2_726, // sfix19_En18 
  input [18:0] Wgt_2_727, // sfix19_En18 
  input [18:0] Wgt_2_728, // sfix19_En18 
  input [18:0] Wgt_2_729, // sfix19_En18 
  input [18:0] Wgt_2_730, // sfix19_En18 
  input [18:0] Wgt_2_731, // sfix19_En18 
  input [18:0] Wgt_2_732, // sfix19_En18 
  input [18:0] Wgt_2_733, // sfix19_En18 
  input [18:0] Wgt_2_734, // sfix19_En18 
  input [18:0] Wgt_2_735, // sfix19_En18 
  input [18:0] Wgt_2_736, // sfix19_En18 
  input [18:0] Wgt_2_737, // sfix19_En18 
  input [18:0] Wgt_2_738, // sfix19_En18 
  input [18:0] Wgt_2_739, // sfix19_En18 
  input [18:0] Wgt_2_740, // sfix19_En18 
  input [18:0] Wgt_2_741, // sfix19_En18 
  input [18:0] Wgt_2_742, // sfix19_En18 
  input [18:0] Wgt_2_743, // sfix19_En18 
  input [18:0] Wgt_2_744, // sfix19_En18 
  input [18:0] Wgt_2_745, // sfix19_En18 
  input [18:0] Wgt_2_746, // sfix19_En18 
  input [18:0] Wgt_2_747, // sfix19_En18 
  input [18:0] Wgt_2_748, // sfix19_En18 
  input [18:0] Wgt_2_749, // sfix19_En18 
  input [18:0] Wgt_2_750, // sfix19_En18 
  input [18:0] Wgt_2_751, // sfix19_En18 
  input [18:0] Wgt_2_752, // sfix19_En18 
  input [18:0] Wgt_2_753, // sfix19_En18 
  input [18:0] Wgt_2_754, // sfix19_En18 
  input [18:0] Wgt_2_755, // sfix19_En18 
  input [18:0] Wgt_2_756, // sfix19_En18 
  input [18:0] Wgt_2_757, // sfix19_En18 
  input [18:0] Wgt_2_758, // sfix19_En18 
  input [18:0] Wgt_2_759, // sfix19_En18 
  input [18:0] Wgt_2_760, // sfix19_En18 
  input [18:0] Wgt_2_761, // sfix19_En18 
  input [18:0] Wgt_2_762, // sfix19_En18 
  input [18:0] Wgt_2_763, // sfix19_En18 
  input [18:0] Wgt_2_764, // sfix19_En18 
  input [18:0] Wgt_2_765, // sfix19_En18 
  input [18:0] Wgt_2_766, // sfix19_En18 
  input [18:0] Wgt_2_767, // sfix19_En18 
  input [18:0] Wgt_2_768, // sfix19_En18 
  input [18:0] Wgt_2_769, // sfix19_En18 
  input [18:0] Wgt_2_770, // sfix19_En18 
  input [18:0] Wgt_2_771, // sfix19_En18 
  input [18:0] Wgt_2_772, // sfix19_En18 
  input [18:0] Wgt_2_773, // sfix19_En18 
  input [18:0] Wgt_2_774, // sfix19_En18 
  input [18:0] Wgt_2_775, // sfix19_En18 
  input [18:0] Wgt_2_776, // sfix19_En18 
  input [18:0] Wgt_2_777, // sfix19_En18 
  input [18:0] Wgt_2_778, // sfix19_En18 
  input [18:0] Wgt_2_779, // sfix19_En18 
  input [18:0] Wgt_2_780, // sfix19_En18 
  input [18:0] Wgt_2_781, // sfix19_En18 
  input [18:0] Wgt_2_782, // sfix19_En18 
  input [18:0] Wgt_2_783, // sfix19_En18 
  input [18:0] Wgt_2_784, // sfix19_En18 
  input [18:0] Wgt_3_0, // sfix19_En18 
  input [18:0] Wgt_3_1, // sfix19_En18 
  input [18:0] Wgt_3_2, // sfix19_En18 
  input [18:0] Wgt_3_3, // sfix19_En18 
  input [18:0] Wgt_3_4, // sfix19_En18 
  input [18:0] Wgt_3_5, // sfix19_En18 
  input [18:0] Wgt_3_6, // sfix19_En18 
  input [18:0] Wgt_3_7, // sfix19_En18 
  input [18:0] Wgt_3_8, // sfix19_En18 
  input [18:0] Wgt_3_9, // sfix19_En18 
  input [18:0] Wgt_3_10, // sfix19_En18 
  input [18:0] Wgt_3_11, // sfix19_En18 
  input [18:0] Wgt_3_12, // sfix19_En18 
  input [18:0] Wgt_3_13, // sfix19_En18 
  input [18:0] Wgt_3_14, // sfix19_En18 
  input [18:0] Wgt_3_15, // sfix19_En18 
  input [18:0] Wgt_3_16, // sfix19_En18 
  input [18:0] Wgt_3_17, // sfix19_En18 
  input [18:0] Wgt_3_18, // sfix19_En18 
  input [18:0] Wgt_3_19, // sfix19_En18 
  input [18:0] Wgt_3_20, // sfix19_En18 
  input [18:0] Wgt_3_21, // sfix19_En18 
  input [18:0] Wgt_3_22, // sfix19_En18 
  input [18:0] Wgt_3_23, // sfix19_En18 
  input [18:0] Wgt_3_24, // sfix19_En18 
  input [18:0] Wgt_3_25, // sfix19_En18 
  input [18:0] Wgt_3_26, // sfix19_En18 
  input [18:0] Wgt_3_27, // sfix19_En18 
  input [18:0] Wgt_3_28, // sfix19_En18 
  input [18:0] Wgt_3_29, // sfix19_En18 
  input [18:0] Wgt_3_30, // sfix19_En18 
  input [18:0] Wgt_3_31, // sfix19_En18 
  input [18:0] Wgt_3_32, // sfix19_En18 
  input [18:0] Wgt_3_33, // sfix19_En18 
  input [18:0] Wgt_3_34, // sfix19_En18 
  input [18:0] Wgt_3_35, // sfix19_En18 
  input [18:0] Wgt_3_36, // sfix19_En18 
  input [18:0] Wgt_3_37, // sfix19_En18 
  input [18:0] Wgt_3_38, // sfix19_En18 
  input [18:0] Wgt_3_39, // sfix19_En18 
  input [18:0] Wgt_3_40, // sfix19_En18 
  input [18:0] Wgt_3_41, // sfix19_En18 
  input [18:0] Wgt_3_42, // sfix19_En18 
  input [18:0] Wgt_3_43, // sfix19_En18 
  input [18:0] Wgt_3_44, // sfix19_En18 
  input [18:0] Wgt_3_45, // sfix19_En18 
  input [18:0] Wgt_3_46, // sfix19_En18 
  input [18:0] Wgt_3_47, // sfix19_En18 
  input [18:0] Wgt_3_48, // sfix19_En18 
  input [18:0] Wgt_3_49, // sfix19_En18 
  input [18:0] Wgt_3_50, // sfix19_En18 
  input [18:0] Wgt_3_51, // sfix19_En18 
  input [18:0] Wgt_3_52, // sfix19_En18 
  input [18:0] Wgt_3_53, // sfix19_En18 
  input [18:0] Wgt_3_54, // sfix19_En18 
  input [18:0] Wgt_3_55, // sfix19_En18 
  input [18:0] Wgt_3_56, // sfix19_En18 
  input [18:0] Wgt_3_57, // sfix19_En18 
  input [18:0] Wgt_3_58, // sfix19_En18 
  input [18:0] Wgt_3_59, // sfix19_En18 
  input [18:0] Wgt_3_60, // sfix19_En18 
  input [18:0] Wgt_3_61, // sfix19_En18 
  input [18:0] Wgt_3_62, // sfix19_En18 
  input [18:0] Wgt_3_63, // sfix19_En18 
  input [18:0] Wgt_3_64, // sfix19_En18 
  input [18:0] Wgt_3_65, // sfix19_En18 
  input [18:0] Wgt_3_66, // sfix19_En18 
  input [18:0] Wgt_3_67, // sfix19_En18 
  input [18:0] Wgt_3_68, // sfix19_En18 
  input [18:0] Wgt_3_69, // sfix19_En18 
  input [18:0] Wgt_3_70, // sfix19_En18 
  input [18:0] Wgt_3_71, // sfix19_En18 
  input [18:0] Wgt_3_72, // sfix19_En18 
  input [18:0] Wgt_3_73, // sfix19_En18 
  input [18:0] Wgt_3_74, // sfix19_En18 
  input [18:0] Wgt_3_75, // sfix19_En18 
  input [18:0] Wgt_3_76, // sfix19_En18 
  input [18:0] Wgt_3_77, // sfix19_En18 
  input [18:0] Wgt_3_78, // sfix19_En18 
  input [18:0] Wgt_3_79, // sfix19_En18 
  input [18:0] Wgt_3_80, // sfix19_En18 
  input [18:0] Wgt_3_81, // sfix19_En18 
  input [18:0] Wgt_3_82, // sfix19_En18 
  input [18:0] Wgt_3_83, // sfix19_En18 
  input [18:0] Wgt_3_84, // sfix19_En18 
  input [18:0] Wgt_3_85, // sfix19_En18 
  input [18:0] Wgt_3_86, // sfix19_En18 
  input [18:0] Wgt_3_87, // sfix19_En18 
  input [18:0] Wgt_3_88, // sfix19_En18 
  input [18:0] Wgt_3_89, // sfix19_En18 
  input [18:0] Wgt_3_90, // sfix19_En18 
  input [18:0] Wgt_3_91, // sfix19_En18 
  input [18:0] Wgt_3_92, // sfix19_En18 
  input [18:0] Wgt_3_93, // sfix19_En18 
  input [18:0] Wgt_3_94, // sfix19_En18 
  input [18:0] Wgt_3_95, // sfix19_En18 
  input [18:0] Wgt_3_96, // sfix19_En18 
  input [18:0] Wgt_3_97, // sfix19_En18 
  input [18:0] Wgt_3_98, // sfix19_En18 
  input [18:0] Wgt_3_99, // sfix19_En18 
  input [18:0] Wgt_3_100, // sfix19_En18 
  input [18:0] Wgt_3_101, // sfix19_En18 
  input [18:0] Wgt_3_102, // sfix19_En18 
  input [18:0] Wgt_3_103, // sfix19_En18 
  input [18:0] Wgt_3_104, // sfix19_En18 
  input [18:0] Wgt_3_105, // sfix19_En18 
  input [18:0] Wgt_3_106, // sfix19_En18 
  input [18:0] Wgt_3_107, // sfix19_En18 
  input [18:0] Wgt_3_108, // sfix19_En18 
  input [18:0] Wgt_3_109, // sfix19_En18 
  input [18:0] Wgt_3_110, // sfix19_En18 
  input [18:0] Wgt_3_111, // sfix19_En18 
  input [18:0] Wgt_3_112, // sfix19_En18 
  input [18:0] Wgt_3_113, // sfix19_En18 
  input [18:0] Wgt_3_114, // sfix19_En18 
  input [18:0] Wgt_3_115, // sfix19_En18 
  input [18:0] Wgt_3_116, // sfix19_En18 
  input [18:0] Wgt_3_117, // sfix19_En18 
  input [18:0] Wgt_3_118, // sfix19_En18 
  input [18:0] Wgt_3_119, // sfix19_En18 
  input [18:0] Wgt_3_120, // sfix19_En18 
  input [18:0] Wgt_3_121, // sfix19_En18 
  input [18:0] Wgt_3_122, // sfix19_En18 
  input [18:0] Wgt_3_123, // sfix19_En18 
  input [18:0] Wgt_3_124, // sfix19_En18 
  input [18:0] Wgt_3_125, // sfix19_En18 
  input [18:0] Wgt_3_126, // sfix19_En18 
  input [18:0] Wgt_3_127, // sfix19_En18 
  input [18:0] Wgt_3_128, // sfix19_En18 
  input [18:0] Wgt_3_129, // sfix19_En18 
  input [18:0] Wgt_3_130, // sfix19_En18 
  input [18:0] Wgt_3_131, // sfix19_En18 
  input [18:0] Wgt_3_132, // sfix19_En18 
  input [18:0] Wgt_3_133, // sfix19_En18 
  input [18:0] Wgt_3_134, // sfix19_En18 
  input [18:0] Wgt_3_135, // sfix19_En18 
  input [18:0] Wgt_3_136, // sfix19_En18 
  input [18:0] Wgt_3_137, // sfix19_En18 
  input [18:0] Wgt_3_138, // sfix19_En18 
  input [18:0] Wgt_3_139, // sfix19_En18 
  input [18:0] Wgt_3_140, // sfix19_En18 
  input [18:0] Wgt_3_141, // sfix19_En18 
  input [18:0] Wgt_3_142, // sfix19_En18 
  input [18:0] Wgt_3_143, // sfix19_En18 
  input [18:0] Wgt_3_144, // sfix19_En18 
  input [18:0] Wgt_3_145, // sfix19_En18 
  input [18:0] Wgt_3_146, // sfix19_En18 
  input [18:0] Wgt_3_147, // sfix19_En18 
  input [18:0] Wgt_3_148, // sfix19_En18 
  input [18:0] Wgt_3_149, // sfix19_En18 
  input [18:0] Wgt_3_150, // sfix19_En18 
  input [18:0] Wgt_3_151, // sfix19_En18 
  input [18:0] Wgt_3_152, // sfix19_En18 
  input [18:0] Wgt_3_153, // sfix19_En18 
  input [18:0] Wgt_3_154, // sfix19_En18 
  input [18:0] Wgt_3_155, // sfix19_En18 
  input [18:0] Wgt_3_156, // sfix19_En18 
  input [18:0] Wgt_3_157, // sfix19_En18 
  input [18:0] Wgt_3_158, // sfix19_En18 
  input [18:0] Wgt_3_159, // sfix19_En18 
  input [18:0] Wgt_3_160, // sfix19_En18 
  input [18:0] Wgt_3_161, // sfix19_En18 
  input [18:0] Wgt_3_162, // sfix19_En18 
  input [18:0] Wgt_3_163, // sfix19_En18 
  input [18:0] Wgt_3_164, // sfix19_En18 
  input [18:0] Wgt_3_165, // sfix19_En18 
  input [18:0] Wgt_3_166, // sfix19_En18 
  input [18:0] Wgt_3_167, // sfix19_En18 
  input [18:0] Wgt_3_168, // sfix19_En18 
  input [18:0] Wgt_3_169, // sfix19_En18 
  input [18:0] Wgt_3_170, // sfix19_En18 
  input [18:0] Wgt_3_171, // sfix19_En18 
  input [18:0] Wgt_3_172, // sfix19_En18 
  input [18:0] Wgt_3_173, // sfix19_En18 
  input [18:0] Wgt_3_174, // sfix19_En18 
  input [18:0] Wgt_3_175, // sfix19_En18 
  input [18:0] Wgt_3_176, // sfix19_En18 
  input [18:0] Wgt_3_177, // sfix19_En18 
  input [18:0] Wgt_3_178, // sfix19_En18 
  input [18:0] Wgt_3_179, // sfix19_En18 
  input [18:0] Wgt_3_180, // sfix19_En18 
  input [18:0] Wgt_3_181, // sfix19_En18 
  input [18:0] Wgt_3_182, // sfix19_En18 
  input [18:0] Wgt_3_183, // sfix19_En18 
  input [18:0] Wgt_3_184, // sfix19_En18 
  input [18:0] Wgt_3_185, // sfix19_En18 
  input [18:0] Wgt_3_186, // sfix19_En18 
  input [18:0] Wgt_3_187, // sfix19_En18 
  input [18:0] Wgt_3_188, // sfix19_En18 
  input [18:0] Wgt_3_189, // sfix19_En18 
  input [18:0] Wgt_3_190, // sfix19_En18 
  input [18:0] Wgt_3_191, // sfix19_En18 
  input [18:0] Wgt_3_192, // sfix19_En18 
  input [18:0] Wgt_3_193, // sfix19_En18 
  input [18:0] Wgt_3_194, // sfix19_En18 
  input [18:0] Wgt_3_195, // sfix19_En18 
  input [18:0] Wgt_3_196, // sfix19_En18 
  input [18:0] Wgt_3_197, // sfix19_En18 
  input [18:0] Wgt_3_198, // sfix19_En18 
  input [18:0] Wgt_3_199, // sfix19_En18 
  input [18:0] Wgt_3_200, // sfix19_En18 
  input [18:0] Wgt_3_201, // sfix19_En18 
  input [18:0] Wgt_3_202, // sfix19_En18 
  input [18:0] Wgt_3_203, // sfix19_En18 
  input [18:0] Wgt_3_204, // sfix19_En18 
  input [18:0] Wgt_3_205, // sfix19_En18 
  input [18:0] Wgt_3_206, // sfix19_En18 
  input [18:0] Wgt_3_207, // sfix19_En18 
  input [18:0] Wgt_3_208, // sfix19_En18 
  input [18:0] Wgt_3_209, // sfix19_En18 
  input [18:0] Wgt_3_210, // sfix19_En18 
  input [18:0] Wgt_3_211, // sfix19_En18 
  input [18:0] Wgt_3_212, // sfix19_En18 
  input [18:0] Wgt_3_213, // sfix19_En18 
  input [18:0] Wgt_3_214, // sfix19_En18 
  input [18:0] Wgt_3_215, // sfix19_En18 
  input [18:0] Wgt_3_216, // sfix19_En18 
  input [18:0] Wgt_3_217, // sfix19_En18 
  input [18:0] Wgt_3_218, // sfix19_En18 
  input [18:0] Wgt_3_219, // sfix19_En18 
  input [18:0] Wgt_3_220, // sfix19_En18 
  input [18:0] Wgt_3_221, // sfix19_En18 
  input [18:0] Wgt_3_222, // sfix19_En18 
  input [18:0] Wgt_3_223, // sfix19_En18 
  input [18:0] Wgt_3_224, // sfix19_En18 
  input [18:0] Wgt_3_225, // sfix19_En18 
  input [18:0] Wgt_3_226, // sfix19_En18 
  input [18:0] Wgt_3_227, // sfix19_En18 
  input [18:0] Wgt_3_228, // sfix19_En18 
  input [18:0] Wgt_3_229, // sfix19_En18 
  input [18:0] Wgt_3_230, // sfix19_En18 
  input [18:0] Wgt_3_231, // sfix19_En18 
  input [18:0] Wgt_3_232, // sfix19_En18 
  input [18:0] Wgt_3_233, // sfix19_En18 
  input [18:0] Wgt_3_234, // sfix19_En18 
  input [18:0] Wgt_3_235, // sfix19_En18 
  input [18:0] Wgt_3_236, // sfix19_En18 
  input [18:0] Wgt_3_237, // sfix19_En18 
  input [18:0] Wgt_3_238, // sfix19_En18 
  input [18:0] Wgt_3_239, // sfix19_En18 
  input [18:0] Wgt_3_240, // sfix19_En18 
  input [18:0] Wgt_3_241, // sfix19_En18 
  input [18:0] Wgt_3_242, // sfix19_En18 
  input [18:0] Wgt_3_243, // sfix19_En18 
  input [18:0] Wgt_3_244, // sfix19_En18 
  input [18:0] Wgt_3_245, // sfix19_En18 
  input [18:0] Wgt_3_246, // sfix19_En18 
  input [18:0] Wgt_3_247, // sfix19_En18 
  input [18:0] Wgt_3_248, // sfix19_En18 
  input [18:0] Wgt_3_249, // sfix19_En18 
  input [18:0] Wgt_3_250, // sfix19_En18 
  input [18:0] Wgt_3_251, // sfix19_En18 
  input [18:0] Wgt_3_252, // sfix19_En18 
  input [18:0] Wgt_3_253, // sfix19_En18 
  input [18:0] Wgt_3_254, // sfix19_En18 
  input [18:0] Wgt_3_255, // sfix19_En18 
  input [18:0] Wgt_3_256, // sfix19_En18 
  input [18:0] Wgt_3_257, // sfix19_En18 
  input [18:0] Wgt_3_258, // sfix19_En18 
  input [18:0] Wgt_3_259, // sfix19_En18 
  input [18:0] Wgt_3_260, // sfix19_En18 
  input [18:0] Wgt_3_261, // sfix19_En18 
  input [18:0] Wgt_3_262, // sfix19_En18 
  input [18:0] Wgt_3_263, // sfix19_En18 
  input [18:0] Wgt_3_264, // sfix19_En18 
  input [18:0] Wgt_3_265, // sfix19_En18 
  input [18:0] Wgt_3_266, // sfix19_En18 
  input [18:0] Wgt_3_267, // sfix19_En18 
  input [18:0] Wgt_3_268, // sfix19_En18 
  input [18:0] Wgt_3_269, // sfix19_En18 
  input [18:0] Wgt_3_270, // sfix19_En18 
  input [18:0] Wgt_3_271, // sfix19_En18 
  input [18:0] Wgt_3_272, // sfix19_En18 
  input [18:0] Wgt_3_273, // sfix19_En18 
  input [18:0] Wgt_3_274, // sfix19_En18 
  input [18:0] Wgt_3_275, // sfix19_En18 
  input [18:0] Wgt_3_276, // sfix19_En18 
  input [18:0] Wgt_3_277, // sfix19_En18 
  input [18:0] Wgt_3_278, // sfix19_En18 
  input [18:0] Wgt_3_279, // sfix19_En18 
  input [18:0] Wgt_3_280, // sfix19_En18 
  input [18:0] Wgt_3_281, // sfix19_En18 
  input [18:0] Wgt_3_282, // sfix19_En18 
  input [18:0] Wgt_3_283, // sfix19_En18 
  input [18:0] Wgt_3_284, // sfix19_En18 
  input [18:0] Wgt_3_285, // sfix19_En18 
  input [18:0] Wgt_3_286, // sfix19_En18 
  input [18:0] Wgt_3_287, // sfix19_En18 
  input [18:0] Wgt_3_288, // sfix19_En18 
  input [18:0] Wgt_3_289, // sfix19_En18 
  input [18:0] Wgt_3_290, // sfix19_En18 
  input [18:0] Wgt_3_291, // sfix19_En18 
  input [18:0] Wgt_3_292, // sfix19_En18 
  input [18:0] Wgt_3_293, // sfix19_En18 
  input [18:0] Wgt_3_294, // sfix19_En18 
  input [18:0] Wgt_3_295, // sfix19_En18 
  input [18:0] Wgt_3_296, // sfix19_En18 
  input [18:0] Wgt_3_297, // sfix19_En18 
  input [18:0] Wgt_3_298, // sfix19_En18 
  input [18:0] Wgt_3_299, // sfix19_En18 
  input [18:0] Wgt_3_300, // sfix19_En18 
  input [18:0] Wgt_3_301, // sfix19_En18 
  input [18:0] Wgt_3_302, // sfix19_En18 
  input [18:0] Wgt_3_303, // sfix19_En18 
  input [18:0] Wgt_3_304, // sfix19_En18 
  input [18:0] Wgt_3_305, // sfix19_En18 
  input [18:0] Wgt_3_306, // sfix19_En18 
  input [18:0] Wgt_3_307, // sfix19_En18 
  input [18:0] Wgt_3_308, // sfix19_En18 
  input [18:0] Wgt_3_309, // sfix19_En18 
  input [18:0] Wgt_3_310, // sfix19_En18 
  input [18:0] Wgt_3_311, // sfix19_En18 
  input [18:0] Wgt_3_312, // sfix19_En18 
  input [18:0] Wgt_3_313, // sfix19_En18 
  input [18:0] Wgt_3_314, // sfix19_En18 
  input [18:0] Wgt_3_315, // sfix19_En18 
  input [18:0] Wgt_3_316, // sfix19_En18 
  input [18:0] Wgt_3_317, // sfix19_En18 
  input [18:0] Wgt_3_318, // sfix19_En18 
  input [18:0] Wgt_3_319, // sfix19_En18 
  input [18:0] Wgt_3_320, // sfix19_En18 
  input [18:0] Wgt_3_321, // sfix19_En18 
  input [18:0] Wgt_3_322, // sfix19_En18 
  input [18:0] Wgt_3_323, // sfix19_En18 
  input [18:0] Wgt_3_324, // sfix19_En18 
  input [18:0] Wgt_3_325, // sfix19_En18 
  input [18:0] Wgt_3_326, // sfix19_En18 
  input [18:0] Wgt_3_327, // sfix19_En18 
  input [18:0] Wgt_3_328, // sfix19_En18 
  input [18:0] Wgt_3_329, // sfix19_En18 
  input [18:0] Wgt_3_330, // sfix19_En18 
  input [18:0] Wgt_3_331, // sfix19_En18 
  input [18:0] Wgt_3_332, // sfix19_En18 
  input [18:0] Wgt_3_333, // sfix19_En18 
  input [18:0] Wgt_3_334, // sfix19_En18 
  input [18:0] Wgt_3_335, // sfix19_En18 
  input [18:0] Wgt_3_336, // sfix19_En18 
  input [18:0] Wgt_3_337, // sfix19_En18 
  input [18:0] Wgt_3_338, // sfix19_En18 
  input [18:0] Wgt_3_339, // sfix19_En18 
  input [18:0] Wgt_3_340, // sfix19_En18 
  input [18:0] Wgt_3_341, // sfix19_En18 
  input [18:0] Wgt_3_342, // sfix19_En18 
  input [18:0] Wgt_3_343, // sfix19_En18 
  input [18:0] Wgt_3_344, // sfix19_En18 
  input [18:0] Wgt_3_345, // sfix19_En18 
  input [18:0] Wgt_3_346, // sfix19_En18 
  input [18:0] Wgt_3_347, // sfix19_En18 
  input [18:0] Wgt_3_348, // sfix19_En18 
  input [18:0] Wgt_3_349, // sfix19_En18 
  input [18:0] Wgt_3_350, // sfix19_En18 
  input [18:0] Wgt_3_351, // sfix19_En18 
  input [18:0] Wgt_3_352, // sfix19_En18 
  input [18:0] Wgt_3_353, // sfix19_En18 
  input [18:0] Wgt_3_354, // sfix19_En18 
  input [18:0] Wgt_3_355, // sfix19_En18 
  input [18:0] Wgt_3_356, // sfix19_En18 
  input [18:0] Wgt_3_357, // sfix19_En18 
  input [18:0] Wgt_3_358, // sfix19_En18 
  input [18:0] Wgt_3_359, // sfix19_En18 
  input [18:0] Wgt_3_360, // sfix19_En18 
  input [18:0] Wgt_3_361, // sfix19_En18 
  input [18:0] Wgt_3_362, // sfix19_En18 
  input [18:0] Wgt_3_363, // sfix19_En18 
  input [18:0] Wgt_3_364, // sfix19_En18 
  input [18:0] Wgt_3_365, // sfix19_En18 
  input [18:0] Wgt_3_366, // sfix19_En18 
  input [18:0] Wgt_3_367, // sfix19_En18 
  input [18:0] Wgt_3_368, // sfix19_En18 
  input [18:0] Wgt_3_369, // sfix19_En18 
  input [18:0] Wgt_3_370, // sfix19_En18 
  input [18:0] Wgt_3_371, // sfix19_En18 
  input [18:0] Wgt_3_372, // sfix19_En18 
  input [18:0] Wgt_3_373, // sfix19_En18 
  input [18:0] Wgt_3_374, // sfix19_En18 
  input [18:0] Wgt_3_375, // sfix19_En18 
  input [18:0] Wgt_3_376, // sfix19_En18 
  input [18:0] Wgt_3_377, // sfix19_En18 
  input [18:0] Wgt_3_378, // sfix19_En18 
  input [18:0] Wgt_3_379, // sfix19_En18 
  input [18:0] Wgt_3_380, // sfix19_En18 
  input [18:0] Wgt_3_381, // sfix19_En18 
  input [18:0] Wgt_3_382, // sfix19_En18 
  input [18:0] Wgt_3_383, // sfix19_En18 
  input [18:0] Wgt_3_384, // sfix19_En18 
  input [18:0] Wgt_3_385, // sfix19_En18 
  input [18:0] Wgt_3_386, // sfix19_En18 
  input [18:0] Wgt_3_387, // sfix19_En18 
  input [18:0] Wgt_3_388, // sfix19_En18 
  input [18:0] Wgt_3_389, // sfix19_En18 
  input [18:0] Wgt_3_390, // sfix19_En18 
  input [18:0] Wgt_3_391, // sfix19_En18 
  input [18:0] Wgt_3_392, // sfix19_En18 
  input [18:0] Wgt_3_393, // sfix19_En18 
  input [18:0] Wgt_3_394, // sfix19_En18 
  input [18:0] Wgt_3_395, // sfix19_En18 
  input [18:0] Wgt_3_396, // sfix19_En18 
  input [18:0] Wgt_3_397, // sfix19_En18 
  input [18:0] Wgt_3_398, // sfix19_En18 
  input [18:0] Wgt_3_399, // sfix19_En18 
  input [18:0] Wgt_3_400, // sfix19_En18 
  input [18:0] Wgt_3_401, // sfix19_En18 
  input [18:0] Wgt_3_402, // sfix19_En18 
  input [18:0] Wgt_3_403, // sfix19_En18 
  input [18:0] Wgt_3_404, // sfix19_En18 
  input [18:0] Wgt_3_405, // sfix19_En18 
  input [18:0] Wgt_3_406, // sfix19_En18 
  input [18:0] Wgt_3_407, // sfix19_En18 
  input [18:0] Wgt_3_408, // sfix19_En18 
  input [18:0] Wgt_3_409, // sfix19_En18 
  input [18:0] Wgt_3_410, // sfix19_En18 
  input [18:0] Wgt_3_411, // sfix19_En18 
  input [18:0] Wgt_3_412, // sfix19_En18 
  input [18:0] Wgt_3_413, // sfix19_En18 
  input [18:0] Wgt_3_414, // sfix19_En18 
  input [18:0] Wgt_3_415, // sfix19_En18 
  input [18:0] Wgt_3_416, // sfix19_En18 
  input [18:0] Wgt_3_417, // sfix19_En18 
  input [18:0] Wgt_3_418, // sfix19_En18 
  input [18:0] Wgt_3_419, // sfix19_En18 
  input [18:0] Wgt_3_420, // sfix19_En18 
  input [18:0] Wgt_3_421, // sfix19_En18 
  input [18:0] Wgt_3_422, // sfix19_En18 
  input [18:0] Wgt_3_423, // sfix19_En18 
  input [18:0] Wgt_3_424, // sfix19_En18 
  input [18:0] Wgt_3_425, // sfix19_En18 
  input [18:0] Wgt_3_426, // sfix19_En18 
  input [18:0] Wgt_3_427, // sfix19_En18 
  input [18:0] Wgt_3_428, // sfix19_En18 
  input [18:0] Wgt_3_429, // sfix19_En18 
  input [18:0] Wgt_3_430, // sfix19_En18 
  input [18:0] Wgt_3_431, // sfix19_En18 
  input [18:0] Wgt_3_432, // sfix19_En18 
  input [18:0] Wgt_3_433, // sfix19_En18 
  input [18:0] Wgt_3_434, // sfix19_En18 
  input [18:0] Wgt_3_435, // sfix19_En18 
  input [18:0] Wgt_3_436, // sfix19_En18 
  input [18:0] Wgt_3_437, // sfix19_En18 
  input [18:0] Wgt_3_438, // sfix19_En18 
  input [18:0] Wgt_3_439, // sfix19_En18 
  input [18:0] Wgt_3_440, // sfix19_En18 
  input [18:0] Wgt_3_441, // sfix19_En18 
  input [18:0] Wgt_3_442, // sfix19_En18 
  input [18:0] Wgt_3_443, // sfix19_En18 
  input [18:0] Wgt_3_444, // sfix19_En18 
  input [18:0] Wgt_3_445, // sfix19_En18 
  input [18:0] Wgt_3_446, // sfix19_En18 
  input [18:0] Wgt_3_447, // sfix19_En18 
  input [18:0] Wgt_3_448, // sfix19_En18 
  input [18:0] Wgt_3_449, // sfix19_En18 
  input [18:0] Wgt_3_450, // sfix19_En18 
  input [18:0] Wgt_3_451, // sfix19_En18 
  input [18:0] Wgt_3_452, // sfix19_En18 
  input [18:0] Wgt_3_453, // sfix19_En18 
  input [18:0] Wgt_3_454, // sfix19_En18 
  input [18:0] Wgt_3_455, // sfix19_En18 
  input [18:0] Wgt_3_456, // sfix19_En18 
  input [18:0] Wgt_3_457, // sfix19_En18 
  input [18:0] Wgt_3_458, // sfix19_En18 
  input [18:0] Wgt_3_459, // sfix19_En18 
  input [18:0] Wgt_3_460, // sfix19_En18 
  input [18:0] Wgt_3_461, // sfix19_En18 
  input [18:0] Wgt_3_462, // sfix19_En18 
  input [18:0] Wgt_3_463, // sfix19_En18 
  input [18:0] Wgt_3_464, // sfix19_En18 
  input [18:0] Wgt_3_465, // sfix19_En18 
  input [18:0] Wgt_3_466, // sfix19_En18 
  input [18:0] Wgt_3_467, // sfix19_En18 
  input [18:0] Wgt_3_468, // sfix19_En18 
  input [18:0] Wgt_3_469, // sfix19_En18 
  input [18:0] Wgt_3_470, // sfix19_En18 
  input [18:0] Wgt_3_471, // sfix19_En18 
  input [18:0] Wgt_3_472, // sfix19_En18 
  input [18:0] Wgt_3_473, // sfix19_En18 
  input [18:0] Wgt_3_474, // sfix19_En18 
  input [18:0] Wgt_3_475, // sfix19_En18 
  input [18:0] Wgt_3_476, // sfix19_En18 
  input [18:0] Wgt_3_477, // sfix19_En18 
  input [18:0] Wgt_3_478, // sfix19_En18 
  input [18:0] Wgt_3_479, // sfix19_En18 
  input [18:0] Wgt_3_480, // sfix19_En18 
  input [18:0] Wgt_3_481, // sfix19_En18 
  input [18:0] Wgt_3_482, // sfix19_En18 
  input [18:0] Wgt_3_483, // sfix19_En18 
  input [18:0] Wgt_3_484, // sfix19_En18 
  input [18:0] Wgt_3_485, // sfix19_En18 
  input [18:0] Wgt_3_486, // sfix19_En18 
  input [18:0] Wgt_3_487, // sfix19_En18 
  input [18:0] Wgt_3_488, // sfix19_En18 
  input [18:0] Wgt_3_489, // sfix19_En18 
  input [18:0] Wgt_3_490, // sfix19_En18 
  input [18:0] Wgt_3_491, // sfix19_En18 
  input [18:0] Wgt_3_492, // sfix19_En18 
  input [18:0] Wgt_3_493, // sfix19_En18 
  input [18:0] Wgt_3_494, // sfix19_En18 
  input [18:0] Wgt_3_495, // sfix19_En18 
  input [18:0] Wgt_3_496, // sfix19_En18 
  input [18:0] Wgt_3_497, // sfix19_En18 
  input [18:0] Wgt_3_498, // sfix19_En18 
  input [18:0] Wgt_3_499, // sfix19_En18 
  input [18:0] Wgt_3_500, // sfix19_En18 
  input [18:0] Wgt_3_501, // sfix19_En18 
  input [18:0] Wgt_3_502, // sfix19_En18 
  input [18:0] Wgt_3_503, // sfix19_En18 
  input [18:0] Wgt_3_504, // sfix19_En18 
  input [18:0] Wgt_3_505, // sfix19_En18 
  input [18:0] Wgt_3_506, // sfix19_En18 
  input [18:0] Wgt_3_507, // sfix19_En18 
  input [18:0] Wgt_3_508, // sfix19_En18 
  input [18:0] Wgt_3_509, // sfix19_En18 
  input [18:0] Wgt_3_510, // sfix19_En18 
  input [18:0] Wgt_3_511, // sfix19_En18 
  input [18:0] Wgt_3_512, // sfix19_En18 
  input [18:0] Wgt_3_513, // sfix19_En18 
  input [18:0] Wgt_3_514, // sfix19_En18 
  input [18:0] Wgt_3_515, // sfix19_En18 
  input [18:0] Wgt_3_516, // sfix19_En18 
  input [18:0] Wgt_3_517, // sfix19_En18 
  input [18:0] Wgt_3_518, // sfix19_En18 
  input [18:0] Wgt_3_519, // sfix19_En18 
  input [18:0] Wgt_3_520, // sfix19_En18 
  input [18:0] Wgt_3_521, // sfix19_En18 
  input [18:0] Wgt_3_522, // sfix19_En18 
  input [18:0] Wgt_3_523, // sfix19_En18 
  input [18:0] Wgt_3_524, // sfix19_En18 
  input [18:0] Wgt_3_525, // sfix19_En18 
  input [18:0] Wgt_3_526, // sfix19_En18 
  input [18:0] Wgt_3_527, // sfix19_En18 
  input [18:0] Wgt_3_528, // sfix19_En18 
  input [18:0] Wgt_3_529, // sfix19_En18 
  input [18:0] Wgt_3_530, // sfix19_En18 
  input [18:0] Wgt_3_531, // sfix19_En18 
  input [18:0] Wgt_3_532, // sfix19_En18 
  input [18:0] Wgt_3_533, // sfix19_En18 
  input [18:0] Wgt_3_534, // sfix19_En18 
  input [18:0] Wgt_3_535, // sfix19_En18 
  input [18:0] Wgt_3_536, // sfix19_En18 
  input [18:0] Wgt_3_537, // sfix19_En18 
  input [18:0] Wgt_3_538, // sfix19_En18 
  input [18:0] Wgt_3_539, // sfix19_En18 
  input [18:0] Wgt_3_540, // sfix19_En18 
  input [18:0] Wgt_3_541, // sfix19_En18 
  input [18:0] Wgt_3_542, // sfix19_En18 
  input [18:0] Wgt_3_543, // sfix19_En18 
  input [18:0] Wgt_3_544, // sfix19_En18 
  input [18:0] Wgt_3_545, // sfix19_En18 
  input [18:0] Wgt_3_546, // sfix19_En18 
  input [18:0] Wgt_3_547, // sfix19_En18 
  input [18:0] Wgt_3_548, // sfix19_En18 
  input [18:0] Wgt_3_549, // sfix19_En18 
  input [18:0] Wgt_3_550, // sfix19_En18 
  input [18:0] Wgt_3_551, // sfix19_En18 
  input [18:0] Wgt_3_552, // sfix19_En18 
  input [18:0] Wgt_3_553, // sfix19_En18 
  input [18:0] Wgt_3_554, // sfix19_En18 
  input [18:0] Wgt_3_555, // sfix19_En18 
  input [18:0] Wgt_3_556, // sfix19_En18 
  input [18:0] Wgt_3_557, // sfix19_En18 
  input [18:0] Wgt_3_558, // sfix19_En18 
  input [18:0] Wgt_3_559, // sfix19_En18 
  input [18:0] Wgt_3_560, // sfix19_En18 
  input [18:0] Wgt_3_561, // sfix19_En18 
  input [18:0] Wgt_3_562, // sfix19_En18 
  input [18:0] Wgt_3_563, // sfix19_En18 
  input [18:0] Wgt_3_564, // sfix19_En18 
  input [18:0] Wgt_3_565, // sfix19_En18 
  input [18:0] Wgt_3_566, // sfix19_En18 
  input [18:0] Wgt_3_567, // sfix19_En18 
  input [18:0] Wgt_3_568, // sfix19_En18 
  input [18:0] Wgt_3_569, // sfix19_En18 
  input [18:0] Wgt_3_570, // sfix19_En18 
  input [18:0] Wgt_3_571, // sfix19_En18 
  input [18:0] Wgt_3_572, // sfix19_En18 
  input [18:0] Wgt_3_573, // sfix19_En18 
  input [18:0] Wgt_3_574, // sfix19_En18 
  input [18:0] Wgt_3_575, // sfix19_En18 
  input [18:0] Wgt_3_576, // sfix19_En18 
  input [18:0] Wgt_3_577, // sfix19_En18 
  input [18:0] Wgt_3_578, // sfix19_En18 
  input [18:0] Wgt_3_579, // sfix19_En18 
  input [18:0] Wgt_3_580, // sfix19_En18 
  input [18:0] Wgt_3_581, // sfix19_En18 
  input [18:0] Wgt_3_582, // sfix19_En18 
  input [18:0] Wgt_3_583, // sfix19_En18 
  input [18:0] Wgt_3_584, // sfix19_En18 
  input [18:0] Wgt_3_585, // sfix19_En18 
  input [18:0] Wgt_3_586, // sfix19_En18 
  input [18:0] Wgt_3_587, // sfix19_En18 
  input [18:0] Wgt_3_588, // sfix19_En18 
  input [18:0] Wgt_3_589, // sfix19_En18 
  input [18:0] Wgt_3_590, // sfix19_En18 
  input [18:0] Wgt_3_591, // sfix19_En18 
  input [18:0] Wgt_3_592, // sfix19_En18 
  input [18:0] Wgt_3_593, // sfix19_En18 
  input [18:0] Wgt_3_594, // sfix19_En18 
  input [18:0] Wgt_3_595, // sfix19_En18 
  input [18:0] Wgt_3_596, // sfix19_En18 
  input [18:0] Wgt_3_597, // sfix19_En18 
  input [18:0] Wgt_3_598, // sfix19_En18 
  input [18:0] Wgt_3_599, // sfix19_En18 
  input [18:0] Wgt_3_600, // sfix19_En18 
  input [18:0] Wgt_3_601, // sfix19_En18 
  input [18:0] Wgt_3_602, // sfix19_En18 
  input [18:0] Wgt_3_603, // sfix19_En18 
  input [18:0] Wgt_3_604, // sfix19_En18 
  input [18:0] Wgt_3_605, // sfix19_En18 
  input [18:0] Wgt_3_606, // sfix19_En18 
  input [18:0] Wgt_3_607, // sfix19_En18 
  input [18:0] Wgt_3_608, // sfix19_En18 
  input [18:0] Wgt_3_609, // sfix19_En18 
  input [18:0] Wgt_3_610, // sfix19_En18 
  input [18:0] Wgt_3_611, // sfix19_En18 
  input [18:0] Wgt_3_612, // sfix19_En18 
  input [18:0] Wgt_3_613, // sfix19_En18 
  input [18:0] Wgt_3_614, // sfix19_En18 
  input [18:0] Wgt_3_615, // sfix19_En18 
  input [18:0] Wgt_3_616, // sfix19_En18 
  input [18:0] Wgt_3_617, // sfix19_En18 
  input [18:0] Wgt_3_618, // sfix19_En18 
  input [18:0] Wgt_3_619, // sfix19_En18 
  input [18:0] Wgt_3_620, // sfix19_En18 
  input [18:0] Wgt_3_621, // sfix19_En18 
  input [18:0] Wgt_3_622, // sfix19_En18 
  input [18:0] Wgt_3_623, // sfix19_En18 
  input [18:0] Wgt_3_624, // sfix19_En18 
  input [18:0] Wgt_3_625, // sfix19_En18 
  input [18:0] Wgt_3_626, // sfix19_En18 
  input [18:0] Wgt_3_627, // sfix19_En18 
  input [18:0] Wgt_3_628, // sfix19_En18 
  input [18:0] Wgt_3_629, // sfix19_En18 
  input [18:0] Wgt_3_630, // sfix19_En18 
  input [18:0] Wgt_3_631, // sfix19_En18 
  input [18:0] Wgt_3_632, // sfix19_En18 
  input [18:0] Wgt_3_633, // sfix19_En18 
  input [18:0] Wgt_3_634, // sfix19_En18 
  input [18:0] Wgt_3_635, // sfix19_En18 
  input [18:0] Wgt_3_636, // sfix19_En18 
  input [18:0] Wgt_3_637, // sfix19_En18 
  input [18:0] Wgt_3_638, // sfix19_En18 
  input [18:0] Wgt_3_639, // sfix19_En18 
  input [18:0] Wgt_3_640, // sfix19_En18 
  input [18:0] Wgt_3_641, // sfix19_En18 
  input [18:0] Wgt_3_642, // sfix19_En18 
  input [18:0] Wgt_3_643, // sfix19_En18 
  input [18:0] Wgt_3_644, // sfix19_En18 
  input [18:0] Wgt_3_645, // sfix19_En18 
  input [18:0] Wgt_3_646, // sfix19_En18 
  input [18:0] Wgt_3_647, // sfix19_En18 
  input [18:0] Wgt_3_648, // sfix19_En18 
  input [18:0] Wgt_3_649, // sfix19_En18 
  input [18:0] Wgt_3_650, // sfix19_En18 
  input [18:0] Wgt_3_651, // sfix19_En18 
  input [18:0] Wgt_3_652, // sfix19_En18 
  input [18:0] Wgt_3_653, // sfix19_En18 
  input [18:0] Wgt_3_654, // sfix19_En18 
  input [18:0] Wgt_3_655, // sfix19_En18 
  input [18:0] Wgt_3_656, // sfix19_En18 
  input [18:0] Wgt_3_657, // sfix19_En18 
  input [18:0] Wgt_3_658, // sfix19_En18 
  input [18:0] Wgt_3_659, // sfix19_En18 
  input [18:0] Wgt_3_660, // sfix19_En18 
  input [18:0] Wgt_3_661, // sfix19_En18 
  input [18:0] Wgt_3_662, // sfix19_En18 
  input [18:0] Wgt_3_663, // sfix19_En18 
  input [18:0] Wgt_3_664, // sfix19_En18 
  input [18:0] Wgt_3_665, // sfix19_En18 
  input [18:0] Wgt_3_666, // sfix19_En18 
  input [18:0] Wgt_3_667, // sfix19_En18 
  input [18:0] Wgt_3_668, // sfix19_En18 
  input [18:0] Wgt_3_669, // sfix19_En18 
  input [18:0] Wgt_3_670, // sfix19_En18 
  input [18:0] Wgt_3_671, // sfix19_En18 
  input [18:0] Wgt_3_672, // sfix19_En18 
  input [18:0] Wgt_3_673, // sfix19_En18 
  input [18:0] Wgt_3_674, // sfix19_En18 
  input [18:0] Wgt_3_675, // sfix19_En18 
  input [18:0] Wgt_3_676, // sfix19_En18 
  input [18:0] Wgt_3_677, // sfix19_En18 
  input [18:0] Wgt_3_678, // sfix19_En18 
  input [18:0] Wgt_3_679, // sfix19_En18 
  input [18:0] Wgt_3_680, // sfix19_En18 
  input [18:0] Wgt_3_681, // sfix19_En18 
  input [18:0] Wgt_3_682, // sfix19_En18 
  input [18:0] Wgt_3_683, // sfix19_En18 
  input [18:0] Wgt_3_684, // sfix19_En18 
  input [18:0] Wgt_3_685, // sfix19_En18 
  input [18:0] Wgt_3_686, // sfix19_En18 
  input [18:0] Wgt_3_687, // sfix19_En18 
  input [18:0] Wgt_3_688, // sfix19_En18 
  input [18:0] Wgt_3_689, // sfix19_En18 
  input [18:0] Wgt_3_690, // sfix19_En18 
  input [18:0] Wgt_3_691, // sfix19_En18 
  input [18:0] Wgt_3_692, // sfix19_En18 
  input [18:0] Wgt_3_693, // sfix19_En18 
  input [18:0] Wgt_3_694, // sfix19_En18 
  input [18:0] Wgt_3_695, // sfix19_En18 
  input [18:0] Wgt_3_696, // sfix19_En18 
  input [18:0] Wgt_3_697, // sfix19_En18 
  input [18:0] Wgt_3_698, // sfix19_En18 
  input [18:0] Wgt_3_699, // sfix19_En18 
  input [18:0] Wgt_3_700, // sfix19_En18 
  input [18:0] Wgt_3_701, // sfix19_En18 
  input [18:0] Wgt_3_702, // sfix19_En18 
  input [18:0] Wgt_3_703, // sfix19_En18 
  input [18:0] Wgt_3_704, // sfix19_En18 
  input [18:0] Wgt_3_705, // sfix19_En18 
  input [18:0] Wgt_3_706, // sfix19_En18 
  input [18:0] Wgt_3_707, // sfix19_En18 
  input [18:0] Wgt_3_708, // sfix19_En18 
  input [18:0] Wgt_3_709, // sfix19_En18 
  input [18:0] Wgt_3_710, // sfix19_En18 
  input [18:0] Wgt_3_711, // sfix19_En18 
  input [18:0] Wgt_3_712, // sfix19_En18 
  input [18:0] Wgt_3_713, // sfix19_En18 
  input [18:0] Wgt_3_714, // sfix19_En18 
  input [18:0] Wgt_3_715, // sfix19_En18 
  input [18:0] Wgt_3_716, // sfix19_En18 
  input [18:0] Wgt_3_717, // sfix19_En18 
  input [18:0] Wgt_3_718, // sfix19_En18 
  input [18:0] Wgt_3_719, // sfix19_En18 
  input [18:0] Wgt_3_720, // sfix19_En18 
  input [18:0] Wgt_3_721, // sfix19_En18 
  input [18:0] Wgt_3_722, // sfix19_En18 
  input [18:0] Wgt_3_723, // sfix19_En18 
  input [18:0] Wgt_3_724, // sfix19_En18 
  input [18:0] Wgt_3_725, // sfix19_En18 
  input [18:0] Wgt_3_726, // sfix19_En18 
  input [18:0] Wgt_3_727, // sfix19_En18 
  input [18:0] Wgt_3_728, // sfix19_En18 
  input [18:0] Wgt_3_729, // sfix19_En18 
  input [18:0] Wgt_3_730, // sfix19_En18 
  input [18:0] Wgt_3_731, // sfix19_En18 
  input [18:0] Wgt_3_732, // sfix19_En18 
  input [18:0] Wgt_3_733, // sfix19_En18 
  input [18:0] Wgt_3_734, // sfix19_En18 
  input [18:0] Wgt_3_735, // sfix19_En18 
  input [18:0] Wgt_3_736, // sfix19_En18 
  input [18:0] Wgt_3_737, // sfix19_En18 
  input [18:0] Wgt_3_738, // sfix19_En18 
  input [18:0] Wgt_3_739, // sfix19_En18 
  input [18:0] Wgt_3_740, // sfix19_En18 
  input [18:0] Wgt_3_741, // sfix19_En18 
  input [18:0] Wgt_3_742, // sfix19_En18 
  input [18:0] Wgt_3_743, // sfix19_En18 
  input [18:0] Wgt_3_744, // sfix19_En18 
  input [18:0] Wgt_3_745, // sfix19_En18 
  input [18:0] Wgt_3_746, // sfix19_En18 
  input [18:0] Wgt_3_747, // sfix19_En18 
  input [18:0] Wgt_3_748, // sfix19_En18 
  input [18:0] Wgt_3_749, // sfix19_En18 
  input [18:0] Wgt_3_750, // sfix19_En18 
  input [18:0] Wgt_3_751, // sfix19_En18 
  input [18:0] Wgt_3_752, // sfix19_En18 
  input [18:0] Wgt_3_753, // sfix19_En18 
  input [18:0] Wgt_3_754, // sfix19_En18 
  input [18:0] Wgt_3_755, // sfix19_En18 
  input [18:0] Wgt_3_756, // sfix19_En18 
  input [18:0] Wgt_3_757, // sfix19_En18 
  input [18:0] Wgt_3_758, // sfix19_En18 
  input [18:0] Wgt_3_759, // sfix19_En18 
  input [18:0] Wgt_3_760, // sfix19_En18 
  input [18:0] Wgt_3_761, // sfix19_En18 
  input [18:0] Wgt_3_762, // sfix19_En18 
  input [18:0] Wgt_3_763, // sfix19_En18 
  input [18:0] Wgt_3_764, // sfix19_En18 
  input [18:0] Wgt_3_765, // sfix19_En18 
  input [18:0] Wgt_3_766, // sfix19_En18 
  input [18:0] Wgt_3_767, // sfix19_En18 
  input [18:0] Wgt_3_768, // sfix19_En18 
  input [18:0] Wgt_3_769, // sfix19_En18 
  input [18:0] Wgt_3_770, // sfix19_En18 
  input [18:0] Wgt_3_771, // sfix19_En18 
  input [18:0] Wgt_3_772, // sfix19_En18 
  input [18:0] Wgt_3_773, // sfix19_En18 
  input [18:0] Wgt_3_774, // sfix19_En18 
  input [18:0] Wgt_3_775, // sfix19_En18 
  input [18:0] Wgt_3_776, // sfix19_En18 
  input [18:0] Wgt_3_777, // sfix19_En18 
  input [18:0] Wgt_3_778, // sfix19_En18 
  input [18:0] Wgt_3_779, // sfix19_En18 
  input [18:0] Wgt_3_780, // sfix19_En18 
  input [18:0] Wgt_3_781, // sfix19_En18 
  input [18:0] Wgt_3_782, // sfix19_En18 
  input [18:0] Wgt_3_783, // sfix19_En18 
  input [18:0] Wgt_3_784, // sfix19_En18 
  input [18:0] Wgt_4_0, // sfix19_En18 
  input [18:0] Wgt_4_1, // sfix19_En18 
  input [18:0] Wgt_4_2, // sfix19_En18 
  input [18:0] Wgt_4_3, // sfix19_En18 
  input [18:0] Wgt_4_4, // sfix19_En18 
  input [18:0] Wgt_4_5, // sfix19_En18 
  input [18:0] Wgt_4_6, // sfix19_En18 
  input [18:0] Wgt_4_7, // sfix19_En18 
  input [18:0] Wgt_4_8, // sfix19_En18 
  input [18:0] Wgt_4_9, // sfix19_En18 
  input [18:0] Wgt_4_10, // sfix19_En18 
  input [18:0] Wgt_4_11, // sfix19_En18 
  input [18:0] Wgt_4_12, // sfix19_En18 
  input [18:0] Wgt_4_13, // sfix19_En18 
  input [18:0] Wgt_4_14, // sfix19_En18 
  input [18:0] Wgt_4_15, // sfix19_En18 
  input [18:0] Wgt_4_16, // sfix19_En18 
  input [18:0] Wgt_4_17, // sfix19_En18 
  input [18:0] Wgt_4_18, // sfix19_En18 
  input [18:0] Wgt_4_19, // sfix19_En18 
  input [18:0] Wgt_4_20, // sfix19_En18 
  input [18:0] Wgt_4_21, // sfix19_En18 
  input [18:0] Wgt_4_22, // sfix19_En18 
  input [18:0] Wgt_4_23, // sfix19_En18 
  input [18:0] Wgt_4_24, // sfix19_En18 
  input [18:0] Wgt_4_25, // sfix19_En18 
  input [18:0] Wgt_4_26, // sfix19_En18 
  input [18:0] Wgt_4_27, // sfix19_En18 
  input [18:0] Wgt_4_28, // sfix19_En18 
  input [18:0] Wgt_4_29, // sfix19_En18 
  input [18:0] Wgt_4_30, // sfix19_En18 
  input [18:0] Wgt_4_31, // sfix19_En18 
  input [18:0] Wgt_4_32, // sfix19_En18 
  input [18:0] Wgt_4_33, // sfix19_En18 
  input [18:0] Wgt_4_34, // sfix19_En18 
  input [18:0] Wgt_4_35, // sfix19_En18 
  input [18:0] Wgt_4_36, // sfix19_En18 
  input [18:0] Wgt_4_37, // sfix19_En18 
  input [18:0] Wgt_4_38, // sfix19_En18 
  input [18:0] Wgt_4_39, // sfix19_En18 
  input [18:0] Wgt_4_40, // sfix19_En18 
  input [18:0] Wgt_4_41, // sfix19_En18 
  input [18:0] Wgt_4_42, // sfix19_En18 
  input [18:0] Wgt_4_43, // sfix19_En18 
  input [18:0] Wgt_4_44, // sfix19_En18 
  input [18:0] Wgt_4_45, // sfix19_En18 
  input [18:0] Wgt_4_46, // sfix19_En18 
  input [18:0] Wgt_4_47, // sfix19_En18 
  input [18:0] Wgt_4_48, // sfix19_En18 
  input [18:0] Wgt_4_49, // sfix19_En18 
  input [18:0] Wgt_4_50, // sfix19_En18 
  input [18:0] Wgt_4_51, // sfix19_En18 
  input [18:0] Wgt_4_52, // sfix19_En18 
  input [18:0] Wgt_4_53, // sfix19_En18 
  input [18:0] Wgt_4_54, // sfix19_En18 
  input [18:0] Wgt_4_55, // sfix19_En18 
  input [18:0] Wgt_4_56, // sfix19_En18 
  input [18:0] Wgt_4_57, // sfix19_En18 
  input [18:0] Wgt_4_58, // sfix19_En18 
  input [18:0] Wgt_4_59, // sfix19_En18 
  input [18:0] Wgt_4_60, // sfix19_En18 
  input [18:0] Wgt_4_61, // sfix19_En18 
  input [18:0] Wgt_4_62, // sfix19_En18 
  input [18:0] Wgt_4_63, // sfix19_En18 
  input [18:0] Wgt_4_64, // sfix19_En18 
  input [18:0] Wgt_4_65, // sfix19_En18 
  input [18:0] Wgt_4_66, // sfix19_En18 
  input [18:0] Wgt_4_67, // sfix19_En18 
  input [18:0] Wgt_4_68, // sfix19_En18 
  input [18:0] Wgt_4_69, // sfix19_En18 
  input [18:0] Wgt_4_70, // sfix19_En18 
  input [18:0] Wgt_4_71, // sfix19_En18 
  input [18:0] Wgt_4_72, // sfix19_En18 
  input [18:0] Wgt_4_73, // sfix19_En18 
  input [18:0] Wgt_4_74, // sfix19_En18 
  input [18:0] Wgt_4_75, // sfix19_En18 
  input [18:0] Wgt_4_76, // sfix19_En18 
  input [18:0] Wgt_4_77, // sfix19_En18 
  input [18:0] Wgt_4_78, // sfix19_En18 
  input [18:0] Wgt_4_79, // sfix19_En18 
  input [18:0] Wgt_4_80, // sfix19_En18 
  input [18:0] Wgt_4_81, // sfix19_En18 
  input [18:0] Wgt_4_82, // sfix19_En18 
  input [18:0] Wgt_4_83, // sfix19_En18 
  input [18:0] Wgt_4_84, // sfix19_En18 
  input [18:0] Wgt_4_85, // sfix19_En18 
  input [18:0] Wgt_4_86, // sfix19_En18 
  input [18:0] Wgt_4_87, // sfix19_En18 
  input [18:0] Wgt_4_88, // sfix19_En18 
  input [18:0] Wgt_4_89, // sfix19_En18 
  input [18:0] Wgt_4_90, // sfix19_En18 
  input [18:0] Wgt_4_91, // sfix19_En18 
  input [18:0] Wgt_4_92, // sfix19_En18 
  input [18:0] Wgt_4_93, // sfix19_En18 
  input [18:0] Wgt_4_94, // sfix19_En18 
  input [18:0] Wgt_4_95, // sfix19_En18 
  input [18:0] Wgt_4_96, // sfix19_En18 
  input [18:0] Wgt_4_97, // sfix19_En18 
  input [18:0] Wgt_4_98, // sfix19_En18 
  input [18:0] Wgt_4_99, // sfix19_En18 
  input [18:0] Wgt_4_100, // sfix19_En18 
  input [18:0] Wgt_4_101, // sfix19_En18 
  input [18:0] Wgt_4_102, // sfix19_En18 
  input [18:0] Wgt_4_103, // sfix19_En18 
  input [18:0] Wgt_4_104, // sfix19_En18 
  input [18:0] Wgt_4_105, // sfix19_En18 
  input [18:0] Wgt_4_106, // sfix19_En18 
  input [18:0] Wgt_4_107, // sfix19_En18 
  input [18:0] Wgt_4_108, // sfix19_En18 
  input [18:0] Wgt_4_109, // sfix19_En18 
  input [18:0] Wgt_4_110, // sfix19_En18 
  input [18:0] Wgt_4_111, // sfix19_En18 
  input [18:0] Wgt_4_112, // sfix19_En18 
  input [18:0] Wgt_4_113, // sfix19_En18 
  input [18:0] Wgt_4_114, // sfix19_En18 
  input [18:0] Wgt_4_115, // sfix19_En18 
  input [18:0] Wgt_4_116, // sfix19_En18 
  input [18:0] Wgt_4_117, // sfix19_En18 
  input [18:0] Wgt_4_118, // sfix19_En18 
  input [18:0] Wgt_4_119, // sfix19_En18 
  input [18:0] Wgt_4_120, // sfix19_En18 
  input [18:0] Wgt_4_121, // sfix19_En18 
  input [18:0] Wgt_4_122, // sfix19_En18 
  input [18:0] Wgt_4_123, // sfix19_En18 
  input [18:0] Wgt_4_124, // sfix19_En18 
  input [18:0] Wgt_4_125, // sfix19_En18 
  input [18:0] Wgt_4_126, // sfix19_En18 
  input [18:0] Wgt_4_127, // sfix19_En18 
  input [18:0] Wgt_4_128, // sfix19_En18 
  input [18:0] Wgt_4_129, // sfix19_En18 
  input [18:0] Wgt_4_130, // sfix19_En18 
  input [18:0] Wgt_4_131, // sfix19_En18 
  input [18:0] Wgt_4_132, // sfix19_En18 
  input [18:0] Wgt_4_133, // sfix19_En18 
  input [18:0] Wgt_4_134, // sfix19_En18 
  input [18:0] Wgt_4_135, // sfix19_En18 
  input [18:0] Wgt_4_136, // sfix19_En18 
  input [18:0] Wgt_4_137, // sfix19_En18 
  input [18:0] Wgt_4_138, // sfix19_En18 
  input [18:0] Wgt_4_139, // sfix19_En18 
  input [18:0] Wgt_4_140, // sfix19_En18 
  input [18:0] Wgt_4_141, // sfix19_En18 
  input [18:0] Wgt_4_142, // sfix19_En18 
  input [18:0] Wgt_4_143, // sfix19_En18 
  input [18:0] Wgt_4_144, // sfix19_En18 
  input [18:0] Wgt_4_145, // sfix19_En18 
  input [18:0] Wgt_4_146, // sfix19_En18 
  input [18:0] Wgt_4_147, // sfix19_En18 
  input [18:0] Wgt_4_148, // sfix19_En18 
  input [18:0] Wgt_4_149, // sfix19_En18 
  input [18:0] Wgt_4_150, // sfix19_En18 
  input [18:0] Wgt_4_151, // sfix19_En18 
  input [18:0] Wgt_4_152, // sfix19_En18 
  input [18:0] Wgt_4_153, // sfix19_En18 
  input [18:0] Wgt_4_154, // sfix19_En18 
  input [18:0] Wgt_4_155, // sfix19_En18 
  input [18:0] Wgt_4_156, // sfix19_En18 
  input [18:0] Wgt_4_157, // sfix19_En18 
  input [18:0] Wgt_4_158, // sfix19_En18 
  input [18:0] Wgt_4_159, // sfix19_En18 
  input [18:0] Wgt_4_160, // sfix19_En18 
  input [18:0] Wgt_4_161, // sfix19_En18 
  input [18:0] Wgt_4_162, // sfix19_En18 
  input [18:0] Wgt_4_163, // sfix19_En18 
  input [18:0] Wgt_4_164, // sfix19_En18 
  input [18:0] Wgt_4_165, // sfix19_En18 
  input [18:0] Wgt_4_166, // sfix19_En18 
  input [18:0] Wgt_4_167, // sfix19_En18 
  input [18:0] Wgt_4_168, // sfix19_En18 
  input [18:0] Wgt_4_169, // sfix19_En18 
  input [18:0] Wgt_4_170, // sfix19_En18 
  input [18:0] Wgt_4_171, // sfix19_En18 
  input [18:0] Wgt_4_172, // sfix19_En18 
  input [18:0] Wgt_4_173, // sfix19_En18 
  input [18:0] Wgt_4_174, // sfix19_En18 
  input [18:0] Wgt_4_175, // sfix19_En18 
  input [18:0] Wgt_4_176, // sfix19_En18 
  input [18:0] Wgt_4_177, // sfix19_En18 
  input [18:0] Wgt_4_178, // sfix19_En18 
  input [18:0] Wgt_4_179, // sfix19_En18 
  input [18:0] Wgt_4_180, // sfix19_En18 
  input [18:0] Wgt_4_181, // sfix19_En18 
  input [18:0] Wgt_4_182, // sfix19_En18 
  input [18:0] Wgt_4_183, // sfix19_En18 
  input [18:0] Wgt_4_184, // sfix19_En18 
  input [18:0] Wgt_4_185, // sfix19_En18 
  input [18:0] Wgt_4_186, // sfix19_En18 
  input [18:0] Wgt_4_187, // sfix19_En18 
  input [18:0] Wgt_4_188, // sfix19_En18 
  input [18:0] Wgt_4_189, // sfix19_En18 
  input [18:0] Wgt_4_190, // sfix19_En18 
  input [18:0] Wgt_4_191, // sfix19_En18 
  input [18:0] Wgt_4_192, // sfix19_En18 
  input [18:0] Wgt_4_193, // sfix19_En18 
  input [18:0] Wgt_4_194, // sfix19_En18 
  input [18:0] Wgt_4_195, // sfix19_En18 
  input [18:0] Wgt_4_196, // sfix19_En18 
  input [18:0] Wgt_4_197, // sfix19_En18 
  input [18:0] Wgt_4_198, // sfix19_En18 
  input [18:0] Wgt_4_199, // sfix19_En18 
  input [18:0] Wgt_4_200, // sfix19_En18 
  input [18:0] Wgt_4_201, // sfix19_En18 
  input [18:0] Wgt_4_202, // sfix19_En18 
  input [18:0] Wgt_4_203, // sfix19_En18 
  input [18:0] Wgt_4_204, // sfix19_En18 
  input [18:0] Wgt_4_205, // sfix19_En18 
  input [18:0] Wgt_4_206, // sfix19_En18 
  input [18:0] Wgt_4_207, // sfix19_En18 
  input [18:0] Wgt_4_208, // sfix19_En18 
  input [18:0] Wgt_4_209, // sfix19_En18 
  input [18:0] Wgt_4_210, // sfix19_En18 
  input [18:0] Wgt_4_211, // sfix19_En18 
  input [18:0] Wgt_4_212, // sfix19_En18 
  input [18:0] Wgt_4_213, // sfix19_En18 
  input [18:0] Wgt_4_214, // sfix19_En18 
  input [18:0] Wgt_4_215, // sfix19_En18 
  input [18:0] Wgt_4_216, // sfix19_En18 
  input [18:0] Wgt_4_217, // sfix19_En18 
  input [18:0] Wgt_4_218, // sfix19_En18 
  input [18:0] Wgt_4_219, // sfix19_En18 
  input [18:0] Wgt_4_220, // sfix19_En18 
  input [18:0] Wgt_4_221, // sfix19_En18 
  input [18:0] Wgt_4_222, // sfix19_En18 
  input [18:0] Wgt_4_223, // sfix19_En18 
  input [18:0] Wgt_4_224, // sfix19_En18 
  input [18:0] Wgt_4_225, // sfix19_En18 
  input [18:0] Wgt_4_226, // sfix19_En18 
  input [18:0] Wgt_4_227, // sfix19_En18 
  input [18:0] Wgt_4_228, // sfix19_En18 
  input [18:0] Wgt_4_229, // sfix19_En18 
  input [18:0] Wgt_4_230, // sfix19_En18 
  input [18:0] Wgt_4_231, // sfix19_En18 
  input [18:0] Wgt_4_232, // sfix19_En18 
  input [18:0] Wgt_4_233, // sfix19_En18 
  input [18:0] Wgt_4_234, // sfix19_En18 
  input [18:0] Wgt_4_235, // sfix19_En18 
  input [18:0] Wgt_4_236, // sfix19_En18 
  input [18:0] Wgt_4_237, // sfix19_En18 
  input [18:0] Wgt_4_238, // sfix19_En18 
  input [18:0] Wgt_4_239, // sfix19_En18 
  input [18:0] Wgt_4_240, // sfix19_En18 
  input [18:0] Wgt_4_241, // sfix19_En18 
  input [18:0] Wgt_4_242, // sfix19_En18 
  input [18:0] Wgt_4_243, // sfix19_En18 
  input [18:0] Wgt_4_244, // sfix19_En18 
  input [18:0] Wgt_4_245, // sfix19_En18 
  input [18:0] Wgt_4_246, // sfix19_En18 
  input [18:0] Wgt_4_247, // sfix19_En18 
  input [18:0] Wgt_4_248, // sfix19_En18 
  input [18:0] Wgt_4_249, // sfix19_En18 
  input [18:0] Wgt_4_250, // sfix19_En18 
  input [18:0] Wgt_4_251, // sfix19_En18 
  input [18:0] Wgt_4_252, // sfix19_En18 
  input [18:0] Wgt_4_253, // sfix19_En18 
  input [18:0] Wgt_4_254, // sfix19_En18 
  input [18:0] Wgt_4_255, // sfix19_En18 
  input [18:0] Wgt_4_256, // sfix19_En18 
  input [18:0] Wgt_4_257, // sfix19_En18 
  input [18:0] Wgt_4_258, // sfix19_En18 
  input [18:0] Wgt_4_259, // sfix19_En18 
  input [18:0] Wgt_4_260, // sfix19_En18 
  input [18:0] Wgt_4_261, // sfix19_En18 
  input [18:0] Wgt_4_262, // sfix19_En18 
  input [18:0] Wgt_4_263, // sfix19_En18 
  input [18:0] Wgt_4_264, // sfix19_En18 
  input [18:0] Wgt_4_265, // sfix19_En18 
  input [18:0] Wgt_4_266, // sfix19_En18 
  input [18:0] Wgt_4_267, // sfix19_En18 
  input [18:0] Wgt_4_268, // sfix19_En18 
  input [18:0] Wgt_4_269, // sfix19_En18 
  input [18:0] Wgt_4_270, // sfix19_En18 
  input [18:0] Wgt_4_271, // sfix19_En18 
  input [18:0] Wgt_4_272, // sfix19_En18 
  input [18:0] Wgt_4_273, // sfix19_En18 
  input [18:0] Wgt_4_274, // sfix19_En18 
  input [18:0] Wgt_4_275, // sfix19_En18 
  input [18:0] Wgt_4_276, // sfix19_En18 
  input [18:0] Wgt_4_277, // sfix19_En18 
  input [18:0] Wgt_4_278, // sfix19_En18 
  input [18:0] Wgt_4_279, // sfix19_En18 
  input [18:0] Wgt_4_280, // sfix19_En18 
  input [18:0] Wgt_4_281, // sfix19_En18 
  input [18:0] Wgt_4_282, // sfix19_En18 
  input [18:0] Wgt_4_283, // sfix19_En18 
  input [18:0] Wgt_4_284, // sfix19_En18 
  input [18:0] Wgt_4_285, // sfix19_En18 
  input [18:0] Wgt_4_286, // sfix19_En18 
  input [18:0] Wgt_4_287, // sfix19_En18 
  input [18:0] Wgt_4_288, // sfix19_En18 
  input [18:0] Wgt_4_289, // sfix19_En18 
  input [18:0] Wgt_4_290, // sfix19_En18 
  input [18:0] Wgt_4_291, // sfix19_En18 
  input [18:0] Wgt_4_292, // sfix19_En18 
  input [18:0] Wgt_4_293, // sfix19_En18 
  input [18:0] Wgt_4_294, // sfix19_En18 
  input [18:0] Wgt_4_295, // sfix19_En18 
  input [18:0] Wgt_4_296, // sfix19_En18 
  input [18:0] Wgt_4_297, // sfix19_En18 
  input [18:0] Wgt_4_298, // sfix19_En18 
  input [18:0] Wgt_4_299, // sfix19_En18 
  input [18:0] Wgt_4_300, // sfix19_En18 
  input [18:0] Wgt_4_301, // sfix19_En18 
  input [18:0] Wgt_4_302, // sfix19_En18 
  input [18:0] Wgt_4_303, // sfix19_En18 
  input [18:0] Wgt_4_304, // sfix19_En18 
  input [18:0] Wgt_4_305, // sfix19_En18 
  input [18:0] Wgt_4_306, // sfix19_En18 
  input [18:0] Wgt_4_307, // sfix19_En18 
  input [18:0] Wgt_4_308, // sfix19_En18 
  input [18:0] Wgt_4_309, // sfix19_En18 
  input [18:0] Wgt_4_310, // sfix19_En18 
  input [18:0] Wgt_4_311, // sfix19_En18 
  input [18:0] Wgt_4_312, // sfix19_En18 
  input [18:0] Wgt_4_313, // sfix19_En18 
  input [18:0] Wgt_4_314, // sfix19_En18 
  input [18:0] Wgt_4_315, // sfix19_En18 
  input [18:0] Wgt_4_316, // sfix19_En18 
  input [18:0] Wgt_4_317, // sfix19_En18 
  input [18:0] Wgt_4_318, // sfix19_En18 
  input [18:0] Wgt_4_319, // sfix19_En18 
  input [18:0] Wgt_4_320, // sfix19_En18 
  input [18:0] Wgt_4_321, // sfix19_En18 
  input [18:0] Wgt_4_322, // sfix19_En18 
  input [18:0] Wgt_4_323, // sfix19_En18 
  input [18:0] Wgt_4_324, // sfix19_En18 
  input [18:0] Wgt_4_325, // sfix19_En18 
  input [18:0] Wgt_4_326, // sfix19_En18 
  input [18:0] Wgt_4_327, // sfix19_En18 
  input [18:0] Wgt_4_328, // sfix19_En18 
  input [18:0] Wgt_4_329, // sfix19_En18 
  input [18:0] Wgt_4_330, // sfix19_En18 
  input [18:0] Wgt_4_331, // sfix19_En18 
  input [18:0] Wgt_4_332, // sfix19_En18 
  input [18:0] Wgt_4_333, // sfix19_En18 
  input [18:0] Wgt_4_334, // sfix19_En18 
  input [18:0] Wgt_4_335, // sfix19_En18 
  input [18:0] Wgt_4_336, // sfix19_En18 
  input [18:0] Wgt_4_337, // sfix19_En18 
  input [18:0] Wgt_4_338, // sfix19_En18 
  input [18:0] Wgt_4_339, // sfix19_En18 
  input [18:0] Wgt_4_340, // sfix19_En18 
  input [18:0] Wgt_4_341, // sfix19_En18 
  input [18:0] Wgt_4_342, // sfix19_En18 
  input [18:0] Wgt_4_343, // sfix19_En18 
  input [18:0] Wgt_4_344, // sfix19_En18 
  input [18:0] Wgt_4_345, // sfix19_En18 
  input [18:0] Wgt_4_346, // sfix19_En18 
  input [18:0] Wgt_4_347, // sfix19_En18 
  input [18:0] Wgt_4_348, // sfix19_En18 
  input [18:0] Wgt_4_349, // sfix19_En18 
  input [18:0] Wgt_4_350, // sfix19_En18 
  input [18:0] Wgt_4_351, // sfix19_En18 
  input [18:0] Wgt_4_352, // sfix19_En18 
  input [18:0] Wgt_4_353, // sfix19_En18 
  input [18:0] Wgt_4_354, // sfix19_En18 
  input [18:0] Wgt_4_355, // sfix19_En18 
  input [18:0] Wgt_4_356, // sfix19_En18 
  input [18:0] Wgt_4_357, // sfix19_En18 
  input [18:0] Wgt_4_358, // sfix19_En18 
  input [18:0] Wgt_4_359, // sfix19_En18 
  input [18:0] Wgt_4_360, // sfix19_En18 
  input [18:0] Wgt_4_361, // sfix19_En18 
  input [18:0] Wgt_4_362, // sfix19_En18 
  input [18:0] Wgt_4_363, // sfix19_En18 
  input [18:0] Wgt_4_364, // sfix19_En18 
  input [18:0] Wgt_4_365, // sfix19_En18 
  input [18:0] Wgt_4_366, // sfix19_En18 
  input [18:0] Wgt_4_367, // sfix19_En18 
  input [18:0] Wgt_4_368, // sfix19_En18 
  input [18:0] Wgt_4_369, // sfix19_En18 
  input [18:0] Wgt_4_370, // sfix19_En18 
  input [18:0] Wgt_4_371, // sfix19_En18 
  input [18:0] Wgt_4_372, // sfix19_En18 
  input [18:0] Wgt_4_373, // sfix19_En18 
  input [18:0] Wgt_4_374, // sfix19_En18 
  input [18:0] Wgt_4_375, // sfix19_En18 
  input [18:0] Wgt_4_376, // sfix19_En18 
  input [18:0] Wgt_4_377, // sfix19_En18 
  input [18:0] Wgt_4_378, // sfix19_En18 
  input [18:0] Wgt_4_379, // sfix19_En18 
  input [18:0] Wgt_4_380, // sfix19_En18 
  input [18:0] Wgt_4_381, // sfix19_En18 
  input [18:0] Wgt_4_382, // sfix19_En18 
  input [18:0] Wgt_4_383, // sfix19_En18 
  input [18:0] Wgt_4_384, // sfix19_En18 
  input [18:0] Wgt_4_385, // sfix19_En18 
  input [18:0] Wgt_4_386, // sfix19_En18 
  input [18:0] Wgt_4_387, // sfix19_En18 
  input [18:0] Wgt_4_388, // sfix19_En18 
  input [18:0] Wgt_4_389, // sfix19_En18 
  input [18:0] Wgt_4_390, // sfix19_En18 
  input [18:0] Wgt_4_391, // sfix19_En18 
  input [18:0] Wgt_4_392, // sfix19_En18 
  input [18:0] Wgt_4_393, // sfix19_En18 
  input [18:0] Wgt_4_394, // sfix19_En18 
  input [18:0] Wgt_4_395, // sfix19_En18 
  input [18:0] Wgt_4_396, // sfix19_En18 
  input [18:0] Wgt_4_397, // sfix19_En18 
  input [18:0] Wgt_4_398, // sfix19_En18 
  input [18:0] Wgt_4_399, // sfix19_En18 
  input [18:0] Wgt_4_400, // sfix19_En18 
  input [18:0] Wgt_4_401, // sfix19_En18 
  input [18:0] Wgt_4_402, // sfix19_En18 
  input [18:0] Wgt_4_403, // sfix19_En18 
  input [18:0] Wgt_4_404, // sfix19_En18 
  input [18:0] Wgt_4_405, // sfix19_En18 
  input [18:0] Wgt_4_406, // sfix19_En18 
  input [18:0] Wgt_4_407, // sfix19_En18 
  input [18:0] Wgt_4_408, // sfix19_En18 
  input [18:0] Wgt_4_409, // sfix19_En18 
  input [18:0] Wgt_4_410, // sfix19_En18 
  input [18:0] Wgt_4_411, // sfix19_En18 
  input [18:0] Wgt_4_412, // sfix19_En18 
  input [18:0] Wgt_4_413, // sfix19_En18 
  input [18:0] Wgt_4_414, // sfix19_En18 
  input [18:0] Wgt_4_415, // sfix19_En18 
  input [18:0] Wgt_4_416, // sfix19_En18 
  input [18:0] Wgt_4_417, // sfix19_En18 
  input [18:0] Wgt_4_418, // sfix19_En18 
  input [18:0] Wgt_4_419, // sfix19_En18 
  input [18:0] Wgt_4_420, // sfix19_En18 
  input [18:0] Wgt_4_421, // sfix19_En18 
  input [18:0] Wgt_4_422, // sfix19_En18 
  input [18:0] Wgt_4_423, // sfix19_En18 
  input [18:0] Wgt_4_424, // sfix19_En18 
  input [18:0] Wgt_4_425, // sfix19_En18 
  input [18:0] Wgt_4_426, // sfix19_En18 
  input [18:0] Wgt_4_427, // sfix19_En18 
  input [18:0] Wgt_4_428, // sfix19_En18 
  input [18:0] Wgt_4_429, // sfix19_En18 
  input [18:0] Wgt_4_430, // sfix19_En18 
  input [18:0] Wgt_4_431, // sfix19_En18 
  input [18:0] Wgt_4_432, // sfix19_En18 
  input [18:0] Wgt_4_433, // sfix19_En18 
  input [18:0] Wgt_4_434, // sfix19_En18 
  input [18:0] Wgt_4_435, // sfix19_En18 
  input [18:0] Wgt_4_436, // sfix19_En18 
  input [18:0] Wgt_4_437, // sfix19_En18 
  input [18:0] Wgt_4_438, // sfix19_En18 
  input [18:0] Wgt_4_439, // sfix19_En18 
  input [18:0] Wgt_4_440, // sfix19_En18 
  input [18:0] Wgt_4_441, // sfix19_En18 
  input [18:0] Wgt_4_442, // sfix19_En18 
  input [18:0] Wgt_4_443, // sfix19_En18 
  input [18:0] Wgt_4_444, // sfix19_En18 
  input [18:0] Wgt_4_445, // sfix19_En18 
  input [18:0] Wgt_4_446, // sfix19_En18 
  input [18:0] Wgt_4_447, // sfix19_En18 
  input [18:0] Wgt_4_448, // sfix19_En18 
  input [18:0] Wgt_4_449, // sfix19_En18 
  input [18:0] Wgt_4_450, // sfix19_En18 
  input [18:0] Wgt_4_451, // sfix19_En18 
  input [18:0] Wgt_4_452, // sfix19_En18 
  input [18:0] Wgt_4_453, // sfix19_En18 
  input [18:0] Wgt_4_454, // sfix19_En18 
  input [18:0] Wgt_4_455, // sfix19_En18 
  input [18:0] Wgt_4_456, // sfix19_En18 
  input [18:0] Wgt_4_457, // sfix19_En18 
  input [18:0] Wgt_4_458, // sfix19_En18 
  input [18:0] Wgt_4_459, // sfix19_En18 
  input [18:0] Wgt_4_460, // sfix19_En18 
  input [18:0] Wgt_4_461, // sfix19_En18 
  input [18:0] Wgt_4_462, // sfix19_En18 
  input [18:0] Wgt_4_463, // sfix19_En18 
  input [18:0] Wgt_4_464, // sfix19_En18 
  input [18:0] Wgt_4_465, // sfix19_En18 
  input [18:0] Wgt_4_466, // sfix19_En18 
  input [18:0] Wgt_4_467, // sfix19_En18 
  input [18:0] Wgt_4_468, // sfix19_En18 
  input [18:0] Wgt_4_469, // sfix19_En18 
  input [18:0] Wgt_4_470, // sfix19_En18 
  input [18:0] Wgt_4_471, // sfix19_En18 
  input [18:0] Wgt_4_472, // sfix19_En18 
  input [18:0] Wgt_4_473, // sfix19_En18 
  input [18:0] Wgt_4_474, // sfix19_En18 
  input [18:0] Wgt_4_475, // sfix19_En18 
  input [18:0] Wgt_4_476, // sfix19_En18 
  input [18:0] Wgt_4_477, // sfix19_En18 
  input [18:0] Wgt_4_478, // sfix19_En18 
  input [18:0] Wgt_4_479, // sfix19_En18 
  input [18:0] Wgt_4_480, // sfix19_En18 
  input [18:0] Wgt_4_481, // sfix19_En18 
  input [18:0] Wgt_4_482, // sfix19_En18 
  input [18:0] Wgt_4_483, // sfix19_En18 
  input [18:0] Wgt_4_484, // sfix19_En18 
  input [18:0] Wgt_4_485, // sfix19_En18 
  input [18:0] Wgt_4_486, // sfix19_En18 
  input [18:0] Wgt_4_487, // sfix19_En18 
  input [18:0] Wgt_4_488, // sfix19_En18 
  input [18:0] Wgt_4_489, // sfix19_En18 
  input [18:0] Wgt_4_490, // sfix19_En18 
  input [18:0] Wgt_4_491, // sfix19_En18 
  input [18:0] Wgt_4_492, // sfix19_En18 
  input [18:0] Wgt_4_493, // sfix19_En18 
  input [18:0] Wgt_4_494, // sfix19_En18 
  input [18:0] Wgt_4_495, // sfix19_En18 
  input [18:0] Wgt_4_496, // sfix19_En18 
  input [18:0] Wgt_4_497, // sfix19_En18 
  input [18:0] Wgt_4_498, // sfix19_En18 
  input [18:0] Wgt_4_499, // sfix19_En18 
  input [18:0] Wgt_4_500, // sfix19_En18 
  input [18:0] Wgt_4_501, // sfix19_En18 
  input [18:0] Wgt_4_502, // sfix19_En18 
  input [18:0] Wgt_4_503, // sfix19_En18 
  input [18:0] Wgt_4_504, // sfix19_En18 
  input [18:0] Wgt_4_505, // sfix19_En18 
  input [18:0] Wgt_4_506, // sfix19_En18 
  input [18:0] Wgt_4_507, // sfix19_En18 
  input [18:0] Wgt_4_508, // sfix19_En18 
  input [18:0] Wgt_4_509, // sfix19_En18 
  input [18:0] Wgt_4_510, // sfix19_En18 
  input [18:0] Wgt_4_511, // sfix19_En18 
  input [18:0] Wgt_4_512, // sfix19_En18 
  input [18:0] Wgt_4_513, // sfix19_En18 
  input [18:0] Wgt_4_514, // sfix19_En18 
  input [18:0] Wgt_4_515, // sfix19_En18 
  input [18:0] Wgt_4_516, // sfix19_En18 
  input [18:0] Wgt_4_517, // sfix19_En18 
  input [18:0] Wgt_4_518, // sfix19_En18 
  input [18:0] Wgt_4_519, // sfix19_En18 
  input [18:0] Wgt_4_520, // sfix19_En18 
  input [18:0] Wgt_4_521, // sfix19_En18 
  input [18:0] Wgt_4_522, // sfix19_En18 
  input [18:0] Wgt_4_523, // sfix19_En18 
  input [18:0] Wgt_4_524, // sfix19_En18 
  input [18:0] Wgt_4_525, // sfix19_En18 
  input [18:0] Wgt_4_526, // sfix19_En18 
  input [18:0] Wgt_4_527, // sfix19_En18 
  input [18:0] Wgt_4_528, // sfix19_En18 
  input [18:0] Wgt_4_529, // sfix19_En18 
  input [18:0] Wgt_4_530, // sfix19_En18 
  input [18:0] Wgt_4_531, // sfix19_En18 
  input [18:0] Wgt_4_532, // sfix19_En18 
  input [18:0] Wgt_4_533, // sfix19_En18 
  input [18:0] Wgt_4_534, // sfix19_En18 
  input [18:0] Wgt_4_535, // sfix19_En18 
  input [18:0] Wgt_4_536, // sfix19_En18 
  input [18:0] Wgt_4_537, // sfix19_En18 
  input [18:0] Wgt_4_538, // sfix19_En18 
  input [18:0] Wgt_4_539, // sfix19_En18 
  input [18:0] Wgt_4_540, // sfix19_En18 
  input [18:0] Wgt_4_541, // sfix19_En18 
  input [18:0] Wgt_4_542, // sfix19_En18 
  input [18:0] Wgt_4_543, // sfix19_En18 
  input [18:0] Wgt_4_544, // sfix19_En18 
  input [18:0] Wgt_4_545, // sfix19_En18 
  input [18:0] Wgt_4_546, // sfix19_En18 
  input [18:0] Wgt_4_547, // sfix19_En18 
  input [18:0] Wgt_4_548, // sfix19_En18 
  input [18:0] Wgt_4_549, // sfix19_En18 
  input [18:0] Wgt_4_550, // sfix19_En18 
  input [18:0] Wgt_4_551, // sfix19_En18 
  input [18:0] Wgt_4_552, // sfix19_En18 
  input [18:0] Wgt_4_553, // sfix19_En18 
  input [18:0] Wgt_4_554, // sfix19_En18 
  input [18:0] Wgt_4_555, // sfix19_En18 
  input [18:0] Wgt_4_556, // sfix19_En18 
  input [18:0] Wgt_4_557, // sfix19_En18 
  input [18:0] Wgt_4_558, // sfix19_En18 
  input [18:0] Wgt_4_559, // sfix19_En18 
  input [18:0] Wgt_4_560, // sfix19_En18 
  input [18:0] Wgt_4_561, // sfix19_En18 
  input [18:0] Wgt_4_562, // sfix19_En18 
  input [18:0] Wgt_4_563, // sfix19_En18 
  input [18:0] Wgt_4_564, // sfix19_En18 
  input [18:0] Wgt_4_565, // sfix19_En18 
  input [18:0] Wgt_4_566, // sfix19_En18 
  input [18:0] Wgt_4_567, // sfix19_En18 
  input [18:0] Wgt_4_568, // sfix19_En18 
  input [18:0] Wgt_4_569, // sfix19_En18 
  input [18:0] Wgt_4_570, // sfix19_En18 
  input [18:0] Wgt_4_571, // sfix19_En18 
  input [18:0] Wgt_4_572, // sfix19_En18 
  input [18:0] Wgt_4_573, // sfix19_En18 
  input [18:0] Wgt_4_574, // sfix19_En18 
  input [18:0] Wgt_4_575, // sfix19_En18 
  input [18:0] Wgt_4_576, // sfix19_En18 
  input [18:0] Wgt_4_577, // sfix19_En18 
  input [18:0] Wgt_4_578, // sfix19_En18 
  input [18:0] Wgt_4_579, // sfix19_En18 
  input [18:0] Wgt_4_580, // sfix19_En18 
  input [18:0] Wgt_4_581, // sfix19_En18 
  input [18:0] Wgt_4_582, // sfix19_En18 
  input [18:0] Wgt_4_583, // sfix19_En18 
  input [18:0] Wgt_4_584, // sfix19_En18 
  input [18:0] Wgt_4_585, // sfix19_En18 
  input [18:0] Wgt_4_586, // sfix19_En18 
  input [18:0] Wgt_4_587, // sfix19_En18 
  input [18:0] Wgt_4_588, // sfix19_En18 
  input [18:0] Wgt_4_589, // sfix19_En18 
  input [18:0] Wgt_4_590, // sfix19_En18 
  input [18:0] Wgt_4_591, // sfix19_En18 
  input [18:0] Wgt_4_592, // sfix19_En18 
  input [18:0] Wgt_4_593, // sfix19_En18 
  input [18:0] Wgt_4_594, // sfix19_En18 
  input [18:0] Wgt_4_595, // sfix19_En18 
  input [18:0] Wgt_4_596, // sfix19_En18 
  input [18:0] Wgt_4_597, // sfix19_En18 
  input [18:0] Wgt_4_598, // sfix19_En18 
  input [18:0] Wgt_4_599, // sfix19_En18 
  input [18:0] Wgt_4_600, // sfix19_En18 
  input [18:0] Wgt_4_601, // sfix19_En18 
  input [18:0] Wgt_4_602, // sfix19_En18 
  input [18:0] Wgt_4_603, // sfix19_En18 
  input [18:0] Wgt_4_604, // sfix19_En18 
  input [18:0] Wgt_4_605, // sfix19_En18 
  input [18:0] Wgt_4_606, // sfix19_En18 
  input [18:0] Wgt_4_607, // sfix19_En18 
  input [18:0] Wgt_4_608, // sfix19_En18 
  input [18:0] Wgt_4_609, // sfix19_En18 
  input [18:0] Wgt_4_610, // sfix19_En18 
  input [18:0] Wgt_4_611, // sfix19_En18 
  input [18:0] Wgt_4_612, // sfix19_En18 
  input [18:0] Wgt_4_613, // sfix19_En18 
  input [18:0] Wgt_4_614, // sfix19_En18 
  input [18:0] Wgt_4_615, // sfix19_En18 
  input [18:0] Wgt_4_616, // sfix19_En18 
  input [18:0] Wgt_4_617, // sfix19_En18 
  input [18:0] Wgt_4_618, // sfix19_En18 
  input [18:0] Wgt_4_619, // sfix19_En18 
  input [18:0] Wgt_4_620, // sfix19_En18 
  input [18:0] Wgt_4_621, // sfix19_En18 
  input [18:0] Wgt_4_622, // sfix19_En18 
  input [18:0] Wgt_4_623, // sfix19_En18 
  input [18:0] Wgt_4_624, // sfix19_En18 
  input [18:0] Wgt_4_625, // sfix19_En18 
  input [18:0] Wgt_4_626, // sfix19_En18 
  input [18:0] Wgt_4_627, // sfix19_En18 
  input [18:0] Wgt_4_628, // sfix19_En18 
  input [18:0] Wgt_4_629, // sfix19_En18 
  input [18:0] Wgt_4_630, // sfix19_En18 
  input [18:0] Wgt_4_631, // sfix19_En18 
  input [18:0] Wgt_4_632, // sfix19_En18 
  input [18:0] Wgt_4_633, // sfix19_En18 
  input [18:0] Wgt_4_634, // sfix19_En18 
  input [18:0] Wgt_4_635, // sfix19_En18 
  input [18:0] Wgt_4_636, // sfix19_En18 
  input [18:0] Wgt_4_637, // sfix19_En18 
  input [18:0] Wgt_4_638, // sfix19_En18 
  input [18:0] Wgt_4_639, // sfix19_En18 
  input [18:0] Wgt_4_640, // sfix19_En18 
  input [18:0] Wgt_4_641, // sfix19_En18 
  input [18:0] Wgt_4_642, // sfix19_En18 
  input [18:0] Wgt_4_643, // sfix19_En18 
  input [18:0] Wgt_4_644, // sfix19_En18 
  input [18:0] Wgt_4_645, // sfix19_En18 
  input [18:0] Wgt_4_646, // sfix19_En18 
  input [18:0] Wgt_4_647, // sfix19_En18 
  input [18:0] Wgt_4_648, // sfix19_En18 
  input [18:0] Wgt_4_649, // sfix19_En18 
  input [18:0] Wgt_4_650, // sfix19_En18 
  input [18:0] Wgt_4_651, // sfix19_En18 
  input [18:0] Wgt_4_652, // sfix19_En18 
  input [18:0] Wgt_4_653, // sfix19_En18 
  input [18:0] Wgt_4_654, // sfix19_En18 
  input [18:0] Wgt_4_655, // sfix19_En18 
  input [18:0] Wgt_4_656, // sfix19_En18 
  input [18:0] Wgt_4_657, // sfix19_En18 
  input [18:0] Wgt_4_658, // sfix19_En18 
  input [18:0] Wgt_4_659, // sfix19_En18 
  input [18:0] Wgt_4_660, // sfix19_En18 
  input [18:0] Wgt_4_661, // sfix19_En18 
  input [18:0] Wgt_4_662, // sfix19_En18 
  input [18:0] Wgt_4_663, // sfix19_En18 
  input [18:0] Wgt_4_664, // sfix19_En18 
  input [18:0] Wgt_4_665, // sfix19_En18 
  input [18:0] Wgt_4_666, // sfix19_En18 
  input [18:0] Wgt_4_667, // sfix19_En18 
  input [18:0] Wgt_4_668, // sfix19_En18 
  input [18:0] Wgt_4_669, // sfix19_En18 
  input [18:0] Wgt_4_670, // sfix19_En18 
  input [18:0] Wgt_4_671, // sfix19_En18 
  input [18:0] Wgt_4_672, // sfix19_En18 
  input [18:0] Wgt_4_673, // sfix19_En18 
  input [18:0] Wgt_4_674, // sfix19_En18 
  input [18:0] Wgt_4_675, // sfix19_En18 
  input [18:0] Wgt_4_676, // sfix19_En18 
  input [18:0] Wgt_4_677, // sfix19_En18 
  input [18:0] Wgt_4_678, // sfix19_En18 
  input [18:0] Wgt_4_679, // sfix19_En18 
  input [18:0] Wgt_4_680, // sfix19_En18 
  input [18:0] Wgt_4_681, // sfix19_En18 
  input [18:0] Wgt_4_682, // sfix19_En18 
  input [18:0] Wgt_4_683, // sfix19_En18 
  input [18:0] Wgt_4_684, // sfix19_En18 
  input [18:0] Wgt_4_685, // sfix19_En18 
  input [18:0] Wgt_4_686, // sfix19_En18 
  input [18:0] Wgt_4_687, // sfix19_En18 
  input [18:0] Wgt_4_688, // sfix19_En18 
  input [18:0] Wgt_4_689, // sfix19_En18 
  input [18:0] Wgt_4_690, // sfix19_En18 
  input [18:0] Wgt_4_691, // sfix19_En18 
  input [18:0] Wgt_4_692, // sfix19_En18 
  input [18:0] Wgt_4_693, // sfix19_En18 
  input [18:0] Wgt_4_694, // sfix19_En18 
  input [18:0] Wgt_4_695, // sfix19_En18 
  input [18:0] Wgt_4_696, // sfix19_En18 
  input [18:0] Wgt_4_697, // sfix19_En18 
  input [18:0] Wgt_4_698, // sfix19_En18 
  input [18:0] Wgt_4_699, // sfix19_En18 
  input [18:0] Wgt_4_700, // sfix19_En18 
  input [18:0] Wgt_4_701, // sfix19_En18 
  input [18:0] Wgt_4_702, // sfix19_En18 
  input [18:0] Wgt_4_703, // sfix19_En18 
  input [18:0] Wgt_4_704, // sfix19_En18 
  input [18:0] Wgt_4_705, // sfix19_En18 
  input [18:0] Wgt_4_706, // sfix19_En18 
  input [18:0] Wgt_4_707, // sfix19_En18 
  input [18:0] Wgt_4_708, // sfix19_En18 
  input [18:0] Wgt_4_709, // sfix19_En18 
  input [18:0] Wgt_4_710, // sfix19_En18 
  input [18:0] Wgt_4_711, // sfix19_En18 
  input [18:0] Wgt_4_712, // sfix19_En18 
  input [18:0] Wgt_4_713, // sfix19_En18 
  input [18:0] Wgt_4_714, // sfix19_En18 
  input [18:0] Wgt_4_715, // sfix19_En18 
  input [18:0] Wgt_4_716, // sfix19_En18 
  input [18:0] Wgt_4_717, // sfix19_En18 
  input [18:0] Wgt_4_718, // sfix19_En18 
  input [18:0] Wgt_4_719, // sfix19_En18 
  input [18:0] Wgt_4_720, // sfix19_En18 
  input [18:0] Wgt_4_721, // sfix19_En18 
  input [18:0] Wgt_4_722, // sfix19_En18 
  input [18:0] Wgt_4_723, // sfix19_En18 
  input [18:0] Wgt_4_724, // sfix19_En18 
  input [18:0] Wgt_4_725, // sfix19_En18 
  input [18:0] Wgt_4_726, // sfix19_En18 
  input [18:0] Wgt_4_727, // sfix19_En18 
  input [18:0] Wgt_4_728, // sfix19_En18 
  input [18:0] Wgt_4_729, // sfix19_En18 
  input [18:0] Wgt_4_730, // sfix19_En18 
  input [18:0] Wgt_4_731, // sfix19_En18 
  input [18:0] Wgt_4_732, // sfix19_En18 
  input [18:0] Wgt_4_733, // sfix19_En18 
  input [18:0] Wgt_4_734, // sfix19_En18 
  input [18:0] Wgt_4_735, // sfix19_En18 
  input [18:0] Wgt_4_736, // sfix19_En18 
  input [18:0] Wgt_4_737, // sfix19_En18 
  input [18:0] Wgt_4_738, // sfix19_En18 
  input [18:0] Wgt_4_739, // sfix19_En18 
  input [18:0] Wgt_4_740, // sfix19_En18 
  input [18:0] Wgt_4_741, // sfix19_En18 
  input [18:0] Wgt_4_742, // sfix19_En18 
  input [18:0] Wgt_4_743, // sfix19_En18 
  input [18:0] Wgt_4_744, // sfix19_En18 
  input [18:0] Wgt_4_745, // sfix19_En18 
  input [18:0] Wgt_4_746, // sfix19_En18 
  input [18:0] Wgt_4_747, // sfix19_En18 
  input [18:0] Wgt_4_748, // sfix19_En18 
  input [18:0] Wgt_4_749, // sfix19_En18 
  input [18:0] Wgt_4_750, // sfix19_En18 
  input [18:0] Wgt_4_751, // sfix19_En18 
  input [18:0] Wgt_4_752, // sfix19_En18 
  input [18:0] Wgt_4_753, // sfix19_En18 
  input [18:0] Wgt_4_754, // sfix19_En18 
  input [18:0] Wgt_4_755, // sfix19_En18 
  input [18:0] Wgt_4_756, // sfix19_En18 
  input [18:0] Wgt_4_757, // sfix19_En18 
  input [18:0] Wgt_4_758, // sfix19_En18 
  input [18:0] Wgt_4_759, // sfix19_En18 
  input [18:0] Wgt_4_760, // sfix19_En18 
  input [18:0] Wgt_4_761, // sfix19_En18 
  input [18:0] Wgt_4_762, // sfix19_En18 
  input [18:0] Wgt_4_763, // sfix19_En18 
  input [18:0] Wgt_4_764, // sfix19_En18 
  input [18:0] Wgt_4_765, // sfix19_En18 
  input [18:0] Wgt_4_766, // sfix19_En18 
  input [18:0] Wgt_4_767, // sfix19_En18 
  input [18:0] Wgt_4_768, // sfix19_En18 
  input [18:0] Wgt_4_769, // sfix19_En18 
  input [18:0] Wgt_4_770, // sfix19_En18 
  input [18:0] Wgt_4_771, // sfix19_En18 
  input [18:0] Wgt_4_772, // sfix19_En18 
  input [18:0] Wgt_4_773, // sfix19_En18 
  input [18:0] Wgt_4_774, // sfix19_En18 
  input [18:0] Wgt_4_775, // sfix19_En18 
  input [18:0] Wgt_4_776, // sfix19_En18 
  input [18:0] Wgt_4_777, // sfix19_En18 
  input [18:0] Wgt_4_778, // sfix19_En18 
  input [18:0] Wgt_4_779, // sfix19_En18 
  input [18:0] Wgt_4_780, // sfix19_En18 
  input [18:0] Wgt_4_781, // sfix19_En18 
  input [18:0] Wgt_4_782, // sfix19_En18 
  input [18:0] Wgt_4_783, // sfix19_En18 
  input [18:0] Wgt_4_784, // sfix19_En18 
  input [18:0] Wgt_5_0, // sfix19_En18 
  input [18:0] Wgt_5_1, // sfix19_En18 
  input [18:0] Wgt_5_2, // sfix19_En18 
  input [18:0] Wgt_5_3, // sfix19_En18 
  input [18:0] Wgt_5_4, // sfix19_En18 
  input [18:0] Wgt_5_5, // sfix19_En18 
  input [18:0] Wgt_5_6, // sfix19_En18 
  input [18:0] Wgt_5_7, // sfix19_En18 
  input [18:0] Wgt_5_8, // sfix19_En18 
  input [18:0] Wgt_5_9, // sfix19_En18 
  input [18:0] Wgt_5_10, // sfix19_En18 
  input [18:0] Wgt_5_11, // sfix19_En18 
  input [18:0] Wgt_5_12, // sfix19_En18 
  input [18:0] Wgt_5_13, // sfix19_En18 
  input [18:0] Wgt_5_14, // sfix19_En18 
  input [18:0] Wgt_5_15, // sfix19_En18 
  input [18:0] Wgt_5_16, // sfix19_En18 
  input [18:0] Wgt_5_17, // sfix19_En18 
  input [18:0] Wgt_5_18, // sfix19_En18 
  input [18:0] Wgt_5_19, // sfix19_En18 
  input [18:0] Wgt_5_20, // sfix19_En18 
  input [18:0] Wgt_5_21, // sfix19_En18 
  input [18:0] Wgt_5_22, // sfix19_En18 
  input [18:0] Wgt_5_23, // sfix19_En18 
  input [18:0] Wgt_5_24, // sfix19_En18 
  input [18:0] Wgt_5_25, // sfix19_En18 
  input [18:0] Wgt_5_26, // sfix19_En18 
  input [18:0] Wgt_5_27, // sfix19_En18 
  input [18:0] Wgt_5_28, // sfix19_En18 
  input [18:0] Wgt_5_29, // sfix19_En18 
  input [18:0] Wgt_5_30, // sfix19_En18 
  input [18:0] Wgt_5_31, // sfix19_En18 
  input [18:0] Wgt_5_32, // sfix19_En18 
  input [18:0] Wgt_5_33, // sfix19_En18 
  input [18:0] Wgt_5_34, // sfix19_En18 
  input [18:0] Wgt_5_35, // sfix19_En18 
  input [18:0] Wgt_5_36, // sfix19_En18 
  input [18:0] Wgt_5_37, // sfix19_En18 
  input [18:0] Wgt_5_38, // sfix19_En18 
  input [18:0] Wgt_5_39, // sfix19_En18 
  input [18:0] Wgt_5_40, // sfix19_En18 
  input [18:0] Wgt_5_41, // sfix19_En18 
  input [18:0] Wgt_5_42, // sfix19_En18 
  input [18:0] Wgt_5_43, // sfix19_En18 
  input [18:0] Wgt_5_44, // sfix19_En18 
  input [18:0] Wgt_5_45, // sfix19_En18 
  input [18:0] Wgt_5_46, // sfix19_En18 
  input [18:0] Wgt_5_47, // sfix19_En18 
  input [18:0] Wgt_5_48, // sfix19_En18 
  input [18:0] Wgt_5_49, // sfix19_En18 
  input [18:0] Wgt_5_50, // sfix19_En18 
  input [18:0] Wgt_5_51, // sfix19_En18 
  input [18:0] Wgt_5_52, // sfix19_En18 
  input [18:0] Wgt_5_53, // sfix19_En18 
  input [18:0] Wgt_5_54, // sfix19_En18 
  input [18:0] Wgt_5_55, // sfix19_En18 
  input [18:0] Wgt_5_56, // sfix19_En18 
  input [18:0] Wgt_5_57, // sfix19_En18 
  input [18:0] Wgt_5_58, // sfix19_En18 
  input [18:0] Wgt_5_59, // sfix19_En18 
  input [18:0] Wgt_5_60, // sfix19_En18 
  input [18:0] Wgt_5_61, // sfix19_En18 
  input [18:0] Wgt_5_62, // sfix19_En18 
  input [18:0] Wgt_5_63, // sfix19_En18 
  input [18:0] Wgt_5_64, // sfix19_En18 
  input [18:0] Wgt_5_65, // sfix19_En18 
  input [18:0] Wgt_5_66, // sfix19_En18 
  input [18:0] Wgt_5_67, // sfix19_En18 
  input [18:0] Wgt_5_68, // sfix19_En18 
  input [18:0] Wgt_5_69, // sfix19_En18 
  input [18:0] Wgt_5_70, // sfix19_En18 
  input [18:0] Wgt_5_71, // sfix19_En18 
  input [18:0] Wgt_5_72, // sfix19_En18 
  input [18:0] Wgt_5_73, // sfix19_En18 
  input [18:0] Wgt_5_74, // sfix19_En18 
  input [18:0] Wgt_5_75, // sfix19_En18 
  input [18:0] Wgt_5_76, // sfix19_En18 
  input [18:0] Wgt_5_77, // sfix19_En18 
  input [18:0] Wgt_5_78, // sfix19_En18 
  input [18:0] Wgt_5_79, // sfix19_En18 
  input [18:0] Wgt_5_80, // sfix19_En18 
  input [18:0] Wgt_5_81, // sfix19_En18 
  input [18:0] Wgt_5_82, // sfix19_En18 
  input [18:0] Wgt_5_83, // sfix19_En18 
  input [18:0] Wgt_5_84, // sfix19_En18 
  input [18:0] Wgt_5_85, // sfix19_En18 
  input [18:0] Wgt_5_86, // sfix19_En18 
  input [18:0] Wgt_5_87, // sfix19_En18 
  input [18:0] Wgt_5_88, // sfix19_En18 
  input [18:0] Wgt_5_89, // sfix19_En18 
  input [18:0] Wgt_5_90, // sfix19_En18 
  input [18:0] Wgt_5_91, // sfix19_En18 
  input [18:0] Wgt_5_92, // sfix19_En18 
  input [18:0] Wgt_5_93, // sfix19_En18 
  input [18:0] Wgt_5_94, // sfix19_En18 
  input [18:0] Wgt_5_95, // sfix19_En18 
  input [18:0] Wgt_5_96, // sfix19_En18 
  input [18:0] Wgt_5_97, // sfix19_En18 
  input [18:0] Wgt_5_98, // sfix19_En18 
  input [18:0] Wgt_5_99, // sfix19_En18 
  input [18:0] Wgt_5_100, // sfix19_En18 
  input [18:0] Wgt_5_101, // sfix19_En18 
  input [18:0] Wgt_5_102, // sfix19_En18 
  input [18:0] Wgt_5_103, // sfix19_En18 
  input [18:0] Wgt_5_104, // sfix19_En18 
  input [18:0] Wgt_5_105, // sfix19_En18 
  input [18:0] Wgt_5_106, // sfix19_En18 
  input [18:0] Wgt_5_107, // sfix19_En18 
  input [18:0] Wgt_5_108, // sfix19_En18 
  input [18:0] Wgt_5_109, // sfix19_En18 
  input [18:0] Wgt_5_110, // sfix19_En18 
  input [18:0] Wgt_5_111, // sfix19_En18 
  input [18:0] Wgt_5_112, // sfix19_En18 
  input [18:0] Wgt_5_113, // sfix19_En18 
  input [18:0] Wgt_5_114, // sfix19_En18 
  input [18:0] Wgt_5_115, // sfix19_En18 
  input [18:0] Wgt_5_116, // sfix19_En18 
  input [18:0] Wgt_5_117, // sfix19_En18 
  input [18:0] Wgt_5_118, // sfix19_En18 
  input [18:0] Wgt_5_119, // sfix19_En18 
  input [18:0] Wgt_5_120, // sfix19_En18 
  input [18:0] Wgt_5_121, // sfix19_En18 
  input [18:0] Wgt_5_122, // sfix19_En18 
  input [18:0] Wgt_5_123, // sfix19_En18 
  input [18:0] Wgt_5_124, // sfix19_En18 
  input [18:0] Wgt_5_125, // sfix19_En18 
  input [18:0] Wgt_5_126, // sfix19_En18 
  input [18:0] Wgt_5_127, // sfix19_En18 
  input [18:0] Wgt_5_128, // sfix19_En18 
  input [18:0] Wgt_5_129, // sfix19_En18 
  input [18:0] Wgt_5_130, // sfix19_En18 
  input [18:0] Wgt_5_131, // sfix19_En18 
  input [18:0] Wgt_5_132, // sfix19_En18 
  input [18:0] Wgt_5_133, // sfix19_En18 
  input [18:0] Wgt_5_134, // sfix19_En18 
  input [18:0] Wgt_5_135, // sfix19_En18 
  input [18:0] Wgt_5_136, // sfix19_En18 
  input [18:0] Wgt_5_137, // sfix19_En18 
  input [18:0] Wgt_5_138, // sfix19_En18 
  input [18:0] Wgt_5_139, // sfix19_En18 
  input [18:0] Wgt_5_140, // sfix19_En18 
  input [18:0] Wgt_5_141, // sfix19_En18 
  input [18:0] Wgt_5_142, // sfix19_En18 
  input [18:0] Wgt_5_143, // sfix19_En18 
  input [18:0] Wgt_5_144, // sfix19_En18 
  input [18:0] Wgt_5_145, // sfix19_En18 
  input [18:0] Wgt_5_146, // sfix19_En18 
  input [18:0] Wgt_5_147, // sfix19_En18 
  input [18:0] Wgt_5_148, // sfix19_En18 
  input [18:0] Wgt_5_149, // sfix19_En18 
  input [18:0] Wgt_5_150, // sfix19_En18 
  input [18:0] Wgt_5_151, // sfix19_En18 
  input [18:0] Wgt_5_152, // sfix19_En18 
  input [18:0] Wgt_5_153, // sfix19_En18 
  input [18:0] Wgt_5_154, // sfix19_En18 
  input [18:0] Wgt_5_155, // sfix19_En18 
  input [18:0] Wgt_5_156, // sfix19_En18 
  input [18:0] Wgt_5_157, // sfix19_En18 
  input [18:0] Wgt_5_158, // sfix19_En18 
  input [18:0] Wgt_5_159, // sfix19_En18 
  input [18:0] Wgt_5_160, // sfix19_En18 
  input [18:0] Wgt_5_161, // sfix19_En18 
  input [18:0] Wgt_5_162, // sfix19_En18 
  input [18:0] Wgt_5_163, // sfix19_En18 
  input [18:0] Wgt_5_164, // sfix19_En18 
  input [18:0] Wgt_5_165, // sfix19_En18 
  input [18:0] Wgt_5_166, // sfix19_En18 
  input [18:0] Wgt_5_167, // sfix19_En18 
  input [18:0] Wgt_5_168, // sfix19_En18 
  input [18:0] Wgt_5_169, // sfix19_En18 
  input [18:0] Wgt_5_170, // sfix19_En18 
  input [18:0] Wgt_5_171, // sfix19_En18 
  input [18:0] Wgt_5_172, // sfix19_En18 
  input [18:0] Wgt_5_173, // sfix19_En18 
  input [18:0] Wgt_5_174, // sfix19_En18 
  input [18:0] Wgt_5_175, // sfix19_En18 
  input [18:0] Wgt_5_176, // sfix19_En18 
  input [18:0] Wgt_5_177, // sfix19_En18 
  input [18:0] Wgt_5_178, // sfix19_En18 
  input [18:0] Wgt_5_179, // sfix19_En18 
  input [18:0] Wgt_5_180, // sfix19_En18 
  input [18:0] Wgt_5_181, // sfix19_En18 
  input [18:0] Wgt_5_182, // sfix19_En18 
  input [18:0] Wgt_5_183, // sfix19_En18 
  input [18:0] Wgt_5_184, // sfix19_En18 
  input [18:0] Wgt_5_185, // sfix19_En18 
  input [18:0] Wgt_5_186, // sfix19_En18 
  input [18:0] Wgt_5_187, // sfix19_En18 
  input [18:0] Wgt_5_188, // sfix19_En18 
  input [18:0] Wgt_5_189, // sfix19_En18 
  input [18:0] Wgt_5_190, // sfix19_En18 
  input [18:0] Wgt_5_191, // sfix19_En18 
  input [18:0] Wgt_5_192, // sfix19_En18 
  input [18:0] Wgt_5_193, // sfix19_En18 
  input [18:0] Wgt_5_194, // sfix19_En18 
  input [18:0] Wgt_5_195, // sfix19_En18 
  input [18:0] Wgt_5_196, // sfix19_En18 
  input [18:0] Wgt_5_197, // sfix19_En18 
  input [18:0] Wgt_5_198, // sfix19_En18 
  input [18:0] Wgt_5_199, // sfix19_En18 
  input [18:0] Wgt_5_200, // sfix19_En18 
  input [18:0] Wgt_5_201, // sfix19_En18 
  input [18:0] Wgt_5_202, // sfix19_En18 
  input [18:0] Wgt_5_203, // sfix19_En18 
  input [18:0] Wgt_5_204, // sfix19_En18 
  input [18:0] Wgt_5_205, // sfix19_En18 
  input [18:0] Wgt_5_206, // sfix19_En18 
  input [18:0] Wgt_5_207, // sfix19_En18 
  input [18:0] Wgt_5_208, // sfix19_En18 
  input [18:0] Wgt_5_209, // sfix19_En18 
  input [18:0] Wgt_5_210, // sfix19_En18 
  input [18:0] Wgt_5_211, // sfix19_En18 
  input [18:0] Wgt_5_212, // sfix19_En18 
  input [18:0] Wgt_5_213, // sfix19_En18 
  input [18:0] Wgt_5_214, // sfix19_En18 
  input [18:0] Wgt_5_215, // sfix19_En18 
  input [18:0] Wgt_5_216, // sfix19_En18 
  input [18:0] Wgt_5_217, // sfix19_En18 
  input [18:0] Wgt_5_218, // sfix19_En18 
  input [18:0] Wgt_5_219, // sfix19_En18 
  input [18:0] Wgt_5_220, // sfix19_En18 
  input [18:0] Wgt_5_221, // sfix19_En18 
  input [18:0] Wgt_5_222, // sfix19_En18 
  input [18:0] Wgt_5_223, // sfix19_En18 
  input [18:0] Wgt_5_224, // sfix19_En18 
  input [18:0] Wgt_5_225, // sfix19_En18 
  input [18:0] Wgt_5_226, // sfix19_En18 
  input [18:0] Wgt_5_227, // sfix19_En18 
  input [18:0] Wgt_5_228, // sfix19_En18 
  input [18:0] Wgt_5_229, // sfix19_En18 
  input [18:0] Wgt_5_230, // sfix19_En18 
  input [18:0] Wgt_5_231, // sfix19_En18 
  input [18:0] Wgt_5_232, // sfix19_En18 
  input [18:0] Wgt_5_233, // sfix19_En18 
  input [18:0] Wgt_5_234, // sfix19_En18 
  input [18:0] Wgt_5_235, // sfix19_En18 
  input [18:0] Wgt_5_236, // sfix19_En18 
  input [18:0] Wgt_5_237, // sfix19_En18 
  input [18:0] Wgt_5_238, // sfix19_En18 
  input [18:0] Wgt_5_239, // sfix19_En18 
  input [18:0] Wgt_5_240, // sfix19_En18 
  input [18:0] Wgt_5_241, // sfix19_En18 
  input [18:0] Wgt_5_242, // sfix19_En18 
  input [18:0] Wgt_5_243, // sfix19_En18 
  input [18:0] Wgt_5_244, // sfix19_En18 
  input [18:0] Wgt_5_245, // sfix19_En18 
  input [18:0] Wgt_5_246, // sfix19_En18 
  input [18:0] Wgt_5_247, // sfix19_En18 
  input [18:0] Wgt_5_248, // sfix19_En18 
  input [18:0] Wgt_5_249, // sfix19_En18 
  input [18:0] Wgt_5_250, // sfix19_En18 
  input [18:0] Wgt_5_251, // sfix19_En18 
  input [18:0] Wgt_5_252, // sfix19_En18 
  input [18:0] Wgt_5_253, // sfix19_En18 
  input [18:0] Wgt_5_254, // sfix19_En18 
  input [18:0] Wgt_5_255, // sfix19_En18 
  input [18:0] Wgt_5_256, // sfix19_En18 
  input [18:0] Wgt_5_257, // sfix19_En18 
  input [18:0] Wgt_5_258, // sfix19_En18 
  input [18:0] Wgt_5_259, // sfix19_En18 
  input [18:0] Wgt_5_260, // sfix19_En18 
  input [18:0] Wgt_5_261, // sfix19_En18 
  input [18:0] Wgt_5_262, // sfix19_En18 
  input [18:0] Wgt_5_263, // sfix19_En18 
  input [18:0] Wgt_5_264, // sfix19_En18 
  input [18:0] Wgt_5_265, // sfix19_En18 
  input [18:0] Wgt_5_266, // sfix19_En18 
  input [18:0] Wgt_5_267, // sfix19_En18 
  input [18:0] Wgt_5_268, // sfix19_En18 
  input [18:0] Wgt_5_269, // sfix19_En18 
  input [18:0] Wgt_5_270, // sfix19_En18 
  input [18:0] Wgt_5_271, // sfix19_En18 
  input [18:0] Wgt_5_272, // sfix19_En18 
  input [18:0] Wgt_5_273, // sfix19_En18 
  input [18:0] Wgt_5_274, // sfix19_En18 
  input [18:0] Wgt_5_275, // sfix19_En18 
  input [18:0] Wgt_5_276, // sfix19_En18 
  input [18:0] Wgt_5_277, // sfix19_En18 
  input [18:0] Wgt_5_278, // sfix19_En18 
  input [18:0] Wgt_5_279, // sfix19_En18 
  input [18:0] Wgt_5_280, // sfix19_En18 
  input [18:0] Wgt_5_281, // sfix19_En18 
  input [18:0] Wgt_5_282, // sfix19_En18 
  input [18:0] Wgt_5_283, // sfix19_En18 
  input [18:0] Wgt_5_284, // sfix19_En18 
  input [18:0] Wgt_5_285, // sfix19_En18 
  input [18:0] Wgt_5_286, // sfix19_En18 
  input [18:0] Wgt_5_287, // sfix19_En18 
  input [18:0] Wgt_5_288, // sfix19_En18 
  input [18:0] Wgt_5_289, // sfix19_En18 
  input [18:0] Wgt_5_290, // sfix19_En18 
  input [18:0] Wgt_5_291, // sfix19_En18 
  input [18:0] Wgt_5_292, // sfix19_En18 
  input [18:0] Wgt_5_293, // sfix19_En18 
  input [18:0] Wgt_5_294, // sfix19_En18 
  input [18:0] Wgt_5_295, // sfix19_En18 
  input [18:0] Wgt_5_296, // sfix19_En18 
  input [18:0] Wgt_5_297, // sfix19_En18 
  input [18:0] Wgt_5_298, // sfix19_En18 
  input [18:0] Wgt_5_299, // sfix19_En18 
  input [18:0] Wgt_5_300, // sfix19_En18 
  input [18:0] Wgt_5_301, // sfix19_En18 
  input [18:0] Wgt_5_302, // sfix19_En18 
  input [18:0] Wgt_5_303, // sfix19_En18 
  input [18:0] Wgt_5_304, // sfix19_En18 
  input [18:0] Wgt_5_305, // sfix19_En18 
  input [18:0] Wgt_5_306, // sfix19_En18 
  input [18:0] Wgt_5_307, // sfix19_En18 
  input [18:0] Wgt_5_308, // sfix19_En18 
  input [18:0] Wgt_5_309, // sfix19_En18 
  input [18:0] Wgt_5_310, // sfix19_En18 
  input [18:0] Wgt_5_311, // sfix19_En18 
  input [18:0] Wgt_5_312, // sfix19_En18 
  input [18:0] Wgt_5_313, // sfix19_En18 
  input [18:0] Wgt_5_314, // sfix19_En18 
  input [18:0] Wgt_5_315, // sfix19_En18 
  input [18:0] Wgt_5_316, // sfix19_En18 
  input [18:0] Wgt_5_317, // sfix19_En18 
  input [18:0] Wgt_5_318, // sfix19_En18 
  input [18:0] Wgt_5_319, // sfix19_En18 
  input [18:0] Wgt_5_320, // sfix19_En18 
  input [18:0] Wgt_5_321, // sfix19_En18 
  input [18:0] Wgt_5_322, // sfix19_En18 
  input [18:0] Wgt_5_323, // sfix19_En18 
  input [18:0] Wgt_5_324, // sfix19_En18 
  input [18:0] Wgt_5_325, // sfix19_En18 
  input [18:0] Wgt_5_326, // sfix19_En18 
  input [18:0] Wgt_5_327, // sfix19_En18 
  input [18:0] Wgt_5_328, // sfix19_En18 
  input [18:0] Wgt_5_329, // sfix19_En18 
  input [18:0] Wgt_5_330, // sfix19_En18 
  input [18:0] Wgt_5_331, // sfix19_En18 
  input [18:0] Wgt_5_332, // sfix19_En18 
  input [18:0] Wgt_5_333, // sfix19_En18 
  input [18:0] Wgt_5_334, // sfix19_En18 
  input [18:0] Wgt_5_335, // sfix19_En18 
  input [18:0] Wgt_5_336, // sfix19_En18 
  input [18:0] Wgt_5_337, // sfix19_En18 
  input [18:0] Wgt_5_338, // sfix19_En18 
  input [18:0] Wgt_5_339, // sfix19_En18 
  input [18:0] Wgt_5_340, // sfix19_En18 
  input [18:0] Wgt_5_341, // sfix19_En18 
  input [18:0] Wgt_5_342, // sfix19_En18 
  input [18:0] Wgt_5_343, // sfix19_En18 
  input [18:0] Wgt_5_344, // sfix19_En18 
  input [18:0] Wgt_5_345, // sfix19_En18 
  input [18:0] Wgt_5_346, // sfix19_En18 
  input [18:0] Wgt_5_347, // sfix19_En18 
  input [18:0] Wgt_5_348, // sfix19_En18 
  input [18:0] Wgt_5_349, // sfix19_En18 
  input [18:0] Wgt_5_350, // sfix19_En18 
  input [18:0] Wgt_5_351, // sfix19_En18 
  input [18:0] Wgt_5_352, // sfix19_En18 
  input [18:0] Wgt_5_353, // sfix19_En18 
  input [18:0] Wgt_5_354, // sfix19_En18 
  input [18:0] Wgt_5_355, // sfix19_En18 
  input [18:0] Wgt_5_356, // sfix19_En18 
  input [18:0] Wgt_5_357, // sfix19_En18 
  input [18:0] Wgt_5_358, // sfix19_En18 
  input [18:0] Wgt_5_359, // sfix19_En18 
  input [18:0] Wgt_5_360, // sfix19_En18 
  input [18:0] Wgt_5_361, // sfix19_En18 
  input [18:0] Wgt_5_362, // sfix19_En18 
  input [18:0] Wgt_5_363, // sfix19_En18 
  input [18:0] Wgt_5_364, // sfix19_En18 
  input [18:0] Wgt_5_365, // sfix19_En18 
  input [18:0] Wgt_5_366, // sfix19_En18 
  input [18:0] Wgt_5_367, // sfix19_En18 
  input [18:0] Wgt_5_368, // sfix19_En18 
  input [18:0] Wgt_5_369, // sfix19_En18 
  input [18:0] Wgt_5_370, // sfix19_En18 
  input [18:0] Wgt_5_371, // sfix19_En18 
  input [18:0] Wgt_5_372, // sfix19_En18 
  input [18:0] Wgt_5_373, // sfix19_En18 
  input [18:0] Wgt_5_374, // sfix19_En18 
  input [18:0] Wgt_5_375, // sfix19_En18 
  input [18:0] Wgt_5_376, // sfix19_En18 
  input [18:0] Wgt_5_377, // sfix19_En18 
  input [18:0] Wgt_5_378, // sfix19_En18 
  input [18:0] Wgt_5_379, // sfix19_En18 
  input [18:0] Wgt_5_380, // sfix19_En18 
  input [18:0] Wgt_5_381, // sfix19_En18 
  input [18:0] Wgt_5_382, // sfix19_En18 
  input [18:0] Wgt_5_383, // sfix19_En18 
  input [18:0] Wgt_5_384, // sfix19_En18 
  input [18:0] Wgt_5_385, // sfix19_En18 
  input [18:0] Wgt_5_386, // sfix19_En18 
  input [18:0] Wgt_5_387, // sfix19_En18 
  input [18:0] Wgt_5_388, // sfix19_En18 
  input [18:0] Wgt_5_389, // sfix19_En18 
  input [18:0] Wgt_5_390, // sfix19_En18 
  input [18:0] Wgt_5_391, // sfix19_En18 
  input [18:0] Wgt_5_392, // sfix19_En18 
  input [18:0] Wgt_5_393, // sfix19_En18 
  input [18:0] Wgt_5_394, // sfix19_En18 
  input [18:0] Wgt_5_395, // sfix19_En18 
  input [18:0] Wgt_5_396, // sfix19_En18 
  input [18:0] Wgt_5_397, // sfix19_En18 
  input [18:0] Wgt_5_398, // sfix19_En18 
  input [18:0] Wgt_5_399, // sfix19_En18 
  input [18:0] Wgt_5_400, // sfix19_En18 
  input [18:0] Wgt_5_401, // sfix19_En18 
  input [18:0] Wgt_5_402, // sfix19_En18 
  input [18:0] Wgt_5_403, // sfix19_En18 
  input [18:0] Wgt_5_404, // sfix19_En18 
  input [18:0] Wgt_5_405, // sfix19_En18 
  input [18:0] Wgt_5_406, // sfix19_En18 
  input [18:0] Wgt_5_407, // sfix19_En18 
  input [18:0] Wgt_5_408, // sfix19_En18 
  input [18:0] Wgt_5_409, // sfix19_En18 
  input [18:0] Wgt_5_410, // sfix19_En18 
  input [18:0] Wgt_5_411, // sfix19_En18 
  input [18:0] Wgt_5_412, // sfix19_En18 
  input [18:0] Wgt_5_413, // sfix19_En18 
  input [18:0] Wgt_5_414, // sfix19_En18 
  input [18:0] Wgt_5_415, // sfix19_En18 
  input [18:0] Wgt_5_416, // sfix19_En18 
  input [18:0] Wgt_5_417, // sfix19_En18 
  input [18:0] Wgt_5_418, // sfix19_En18 
  input [18:0] Wgt_5_419, // sfix19_En18 
  input [18:0] Wgt_5_420, // sfix19_En18 
  input [18:0] Wgt_5_421, // sfix19_En18 
  input [18:0] Wgt_5_422, // sfix19_En18 
  input [18:0] Wgt_5_423, // sfix19_En18 
  input [18:0] Wgt_5_424, // sfix19_En18 
  input [18:0] Wgt_5_425, // sfix19_En18 
  input [18:0] Wgt_5_426, // sfix19_En18 
  input [18:0] Wgt_5_427, // sfix19_En18 
  input [18:0] Wgt_5_428, // sfix19_En18 
  input [18:0] Wgt_5_429, // sfix19_En18 
  input [18:0] Wgt_5_430, // sfix19_En18 
  input [18:0] Wgt_5_431, // sfix19_En18 
  input [18:0] Wgt_5_432, // sfix19_En18 
  input [18:0] Wgt_5_433, // sfix19_En18 
  input [18:0] Wgt_5_434, // sfix19_En18 
  input [18:0] Wgt_5_435, // sfix19_En18 
  input [18:0] Wgt_5_436, // sfix19_En18 
  input [18:0] Wgt_5_437, // sfix19_En18 
  input [18:0] Wgt_5_438, // sfix19_En18 
  input [18:0] Wgt_5_439, // sfix19_En18 
  input [18:0] Wgt_5_440, // sfix19_En18 
  input [18:0] Wgt_5_441, // sfix19_En18 
  input [18:0] Wgt_5_442, // sfix19_En18 
  input [18:0] Wgt_5_443, // sfix19_En18 
  input [18:0] Wgt_5_444, // sfix19_En18 
  input [18:0] Wgt_5_445, // sfix19_En18 
  input [18:0] Wgt_5_446, // sfix19_En18 
  input [18:0] Wgt_5_447, // sfix19_En18 
  input [18:0] Wgt_5_448, // sfix19_En18 
  input [18:0] Wgt_5_449, // sfix19_En18 
  input [18:0] Wgt_5_450, // sfix19_En18 
  input [18:0] Wgt_5_451, // sfix19_En18 
  input [18:0] Wgt_5_452, // sfix19_En18 
  input [18:0] Wgt_5_453, // sfix19_En18 
  input [18:0] Wgt_5_454, // sfix19_En18 
  input [18:0] Wgt_5_455, // sfix19_En18 
  input [18:0] Wgt_5_456, // sfix19_En18 
  input [18:0] Wgt_5_457, // sfix19_En18 
  input [18:0] Wgt_5_458, // sfix19_En18 
  input [18:0] Wgt_5_459, // sfix19_En18 
  input [18:0] Wgt_5_460, // sfix19_En18 
  input [18:0] Wgt_5_461, // sfix19_En18 
  input [18:0] Wgt_5_462, // sfix19_En18 
  input [18:0] Wgt_5_463, // sfix19_En18 
  input [18:0] Wgt_5_464, // sfix19_En18 
  input [18:0] Wgt_5_465, // sfix19_En18 
  input [18:0] Wgt_5_466, // sfix19_En18 
  input [18:0] Wgt_5_467, // sfix19_En18 
  input [18:0] Wgt_5_468, // sfix19_En18 
  input [18:0] Wgt_5_469, // sfix19_En18 
  input [18:0] Wgt_5_470, // sfix19_En18 
  input [18:0] Wgt_5_471, // sfix19_En18 
  input [18:0] Wgt_5_472, // sfix19_En18 
  input [18:0] Wgt_5_473, // sfix19_En18 
  input [18:0] Wgt_5_474, // sfix19_En18 
  input [18:0] Wgt_5_475, // sfix19_En18 
  input [18:0] Wgt_5_476, // sfix19_En18 
  input [18:0] Wgt_5_477, // sfix19_En18 
  input [18:0] Wgt_5_478, // sfix19_En18 
  input [18:0] Wgt_5_479, // sfix19_En18 
  input [18:0] Wgt_5_480, // sfix19_En18 
  input [18:0] Wgt_5_481, // sfix19_En18 
  input [18:0] Wgt_5_482, // sfix19_En18 
  input [18:0] Wgt_5_483, // sfix19_En18 
  input [18:0] Wgt_5_484, // sfix19_En18 
  input [18:0] Wgt_5_485, // sfix19_En18 
  input [18:0] Wgt_5_486, // sfix19_En18 
  input [18:0] Wgt_5_487, // sfix19_En18 
  input [18:0] Wgt_5_488, // sfix19_En18 
  input [18:0] Wgt_5_489, // sfix19_En18 
  input [18:0] Wgt_5_490, // sfix19_En18 
  input [18:0] Wgt_5_491, // sfix19_En18 
  input [18:0] Wgt_5_492, // sfix19_En18 
  input [18:0] Wgt_5_493, // sfix19_En18 
  input [18:0] Wgt_5_494, // sfix19_En18 
  input [18:0] Wgt_5_495, // sfix19_En18 
  input [18:0] Wgt_5_496, // sfix19_En18 
  input [18:0] Wgt_5_497, // sfix19_En18 
  input [18:0] Wgt_5_498, // sfix19_En18 
  input [18:0] Wgt_5_499, // sfix19_En18 
  input [18:0] Wgt_5_500, // sfix19_En18 
  input [18:0] Wgt_5_501, // sfix19_En18 
  input [18:0] Wgt_5_502, // sfix19_En18 
  input [18:0] Wgt_5_503, // sfix19_En18 
  input [18:0] Wgt_5_504, // sfix19_En18 
  input [18:0] Wgt_5_505, // sfix19_En18 
  input [18:0] Wgt_5_506, // sfix19_En18 
  input [18:0] Wgt_5_507, // sfix19_En18 
  input [18:0] Wgt_5_508, // sfix19_En18 
  input [18:0] Wgt_5_509, // sfix19_En18 
  input [18:0] Wgt_5_510, // sfix19_En18 
  input [18:0] Wgt_5_511, // sfix19_En18 
  input [18:0] Wgt_5_512, // sfix19_En18 
  input [18:0] Wgt_5_513, // sfix19_En18 
  input [18:0] Wgt_5_514, // sfix19_En18 
  input [18:0] Wgt_5_515, // sfix19_En18 
  input [18:0] Wgt_5_516, // sfix19_En18 
  input [18:0] Wgt_5_517, // sfix19_En18 
  input [18:0] Wgt_5_518, // sfix19_En18 
  input [18:0] Wgt_5_519, // sfix19_En18 
  input [18:0] Wgt_5_520, // sfix19_En18 
  input [18:0] Wgt_5_521, // sfix19_En18 
  input [18:0] Wgt_5_522, // sfix19_En18 
  input [18:0] Wgt_5_523, // sfix19_En18 
  input [18:0] Wgt_5_524, // sfix19_En18 
  input [18:0] Wgt_5_525, // sfix19_En18 
  input [18:0] Wgt_5_526, // sfix19_En18 
  input [18:0] Wgt_5_527, // sfix19_En18 
  input [18:0] Wgt_5_528, // sfix19_En18 
  input [18:0] Wgt_5_529, // sfix19_En18 
  input [18:0] Wgt_5_530, // sfix19_En18 
  input [18:0] Wgt_5_531, // sfix19_En18 
  input [18:0] Wgt_5_532, // sfix19_En18 
  input [18:0] Wgt_5_533, // sfix19_En18 
  input [18:0] Wgt_5_534, // sfix19_En18 
  input [18:0] Wgt_5_535, // sfix19_En18 
  input [18:0] Wgt_5_536, // sfix19_En18 
  input [18:0] Wgt_5_537, // sfix19_En18 
  input [18:0] Wgt_5_538, // sfix19_En18 
  input [18:0] Wgt_5_539, // sfix19_En18 
  input [18:0] Wgt_5_540, // sfix19_En18 
  input [18:0] Wgt_5_541, // sfix19_En18 
  input [18:0] Wgt_5_542, // sfix19_En18 
  input [18:0] Wgt_5_543, // sfix19_En18 
  input [18:0] Wgt_5_544, // sfix19_En18 
  input [18:0] Wgt_5_545, // sfix19_En18 
  input [18:0] Wgt_5_546, // sfix19_En18 
  input [18:0] Wgt_5_547, // sfix19_En18 
  input [18:0] Wgt_5_548, // sfix19_En18 
  input [18:0] Wgt_5_549, // sfix19_En18 
  input [18:0] Wgt_5_550, // sfix19_En18 
  input [18:0] Wgt_5_551, // sfix19_En18 
  input [18:0] Wgt_5_552, // sfix19_En18 
  input [18:0] Wgt_5_553, // sfix19_En18 
  input [18:0] Wgt_5_554, // sfix19_En18 
  input [18:0] Wgt_5_555, // sfix19_En18 
  input [18:0] Wgt_5_556, // sfix19_En18 
  input [18:0] Wgt_5_557, // sfix19_En18 
  input [18:0] Wgt_5_558, // sfix19_En18 
  input [18:0] Wgt_5_559, // sfix19_En18 
  input [18:0] Wgt_5_560, // sfix19_En18 
  input [18:0] Wgt_5_561, // sfix19_En18 
  input [18:0] Wgt_5_562, // sfix19_En18 
  input [18:0] Wgt_5_563, // sfix19_En18 
  input [18:0] Wgt_5_564, // sfix19_En18 
  input [18:0] Wgt_5_565, // sfix19_En18 
  input [18:0] Wgt_5_566, // sfix19_En18 
  input [18:0] Wgt_5_567, // sfix19_En18 
  input [18:0] Wgt_5_568, // sfix19_En18 
  input [18:0] Wgt_5_569, // sfix19_En18 
  input [18:0] Wgt_5_570, // sfix19_En18 
  input [18:0] Wgt_5_571, // sfix19_En18 
  input [18:0] Wgt_5_572, // sfix19_En18 
  input [18:0] Wgt_5_573, // sfix19_En18 
  input [18:0] Wgt_5_574, // sfix19_En18 
  input [18:0] Wgt_5_575, // sfix19_En18 
  input [18:0] Wgt_5_576, // sfix19_En18 
  input [18:0] Wgt_5_577, // sfix19_En18 
  input [18:0] Wgt_5_578, // sfix19_En18 
  input [18:0] Wgt_5_579, // sfix19_En18 
  input [18:0] Wgt_5_580, // sfix19_En18 
  input [18:0] Wgt_5_581, // sfix19_En18 
  input [18:0] Wgt_5_582, // sfix19_En18 
  input [18:0] Wgt_5_583, // sfix19_En18 
  input [18:0] Wgt_5_584, // sfix19_En18 
  input [18:0] Wgt_5_585, // sfix19_En18 
  input [18:0] Wgt_5_586, // sfix19_En18 
  input [18:0] Wgt_5_587, // sfix19_En18 
  input [18:0] Wgt_5_588, // sfix19_En18 
  input [18:0] Wgt_5_589, // sfix19_En18 
  input [18:0] Wgt_5_590, // sfix19_En18 
  input [18:0] Wgt_5_591, // sfix19_En18 
  input [18:0] Wgt_5_592, // sfix19_En18 
  input [18:0] Wgt_5_593, // sfix19_En18 
  input [18:0] Wgt_5_594, // sfix19_En18 
  input [18:0] Wgt_5_595, // sfix19_En18 
  input [18:0] Wgt_5_596, // sfix19_En18 
  input [18:0] Wgt_5_597, // sfix19_En18 
  input [18:0] Wgt_5_598, // sfix19_En18 
  input [18:0] Wgt_5_599, // sfix19_En18 
  input [18:0] Wgt_5_600, // sfix19_En18 
  input [18:0] Wgt_5_601, // sfix19_En18 
  input [18:0] Wgt_5_602, // sfix19_En18 
  input [18:0] Wgt_5_603, // sfix19_En18 
  input [18:0] Wgt_5_604, // sfix19_En18 
  input [18:0] Wgt_5_605, // sfix19_En18 
  input [18:0] Wgt_5_606, // sfix19_En18 
  input [18:0] Wgt_5_607, // sfix19_En18 
  input [18:0] Wgt_5_608, // sfix19_En18 
  input [18:0] Wgt_5_609, // sfix19_En18 
  input [18:0] Wgt_5_610, // sfix19_En18 
  input [18:0] Wgt_5_611, // sfix19_En18 
  input [18:0] Wgt_5_612, // sfix19_En18 
  input [18:0] Wgt_5_613, // sfix19_En18 
  input [18:0] Wgt_5_614, // sfix19_En18 
  input [18:0] Wgt_5_615, // sfix19_En18 
  input [18:0] Wgt_5_616, // sfix19_En18 
  input [18:0] Wgt_5_617, // sfix19_En18 
  input [18:0] Wgt_5_618, // sfix19_En18 
  input [18:0] Wgt_5_619, // sfix19_En18 
  input [18:0] Wgt_5_620, // sfix19_En18 
  input [18:0] Wgt_5_621, // sfix19_En18 
  input [18:0] Wgt_5_622, // sfix19_En18 
  input [18:0] Wgt_5_623, // sfix19_En18 
  input [18:0] Wgt_5_624, // sfix19_En18 
  input [18:0] Wgt_5_625, // sfix19_En18 
  input [18:0] Wgt_5_626, // sfix19_En18 
  input [18:0] Wgt_5_627, // sfix19_En18 
  input [18:0] Wgt_5_628, // sfix19_En18 
  input [18:0] Wgt_5_629, // sfix19_En18 
  input [18:0] Wgt_5_630, // sfix19_En18 
  input [18:0] Wgt_5_631, // sfix19_En18 
  input [18:0] Wgt_5_632, // sfix19_En18 
  input [18:0] Wgt_5_633, // sfix19_En18 
  input [18:0] Wgt_5_634, // sfix19_En18 
  input [18:0] Wgt_5_635, // sfix19_En18 
  input [18:0] Wgt_5_636, // sfix19_En18 
  input [18:0] Wgt_5_637, // sfix19_En18 
  input [18:0] Wgt_5_638, // sfix19_En18 
  input [18:0] Wgt_5_639, // sfix19_En18 
  input [18:0] Wgt_5_640, // sfix19_En18 
  input [18:0] Wgt_5_641, // sfix19_En18 
  input [18:0] Wgt_5_642, // sfix19_En18 
  input [18:0] Wgt_5_643, // sfix19_En18 
  input [18:0] Wgt_5_644, // sfix19_En18 
  input [18:0] Wgt_5_645, // sfix19_En18 
  input [18:0] Wgt_5_646, // sfix19_En18 
  input [18:0] Wgt_5_647, // sfix19_En18 
  input [18:0] Wgt_5_648, // sfix19_En18 
  input [18:0] Wgt_5_649, // sfix19_En18 
  input [18:0] Wgt_5_650, // sfix19_En18 
  input [18:0] Wgt_5_651, // sfix19_En18 
  input [18:0] Wgt_5_652, // sfix19_En18 
  input [18:0] Wgt_5_653, // sfix19_En18 
  input [18:0] Wgt_5_654, // sfix19_En18 
  input [18:0] Wgt_5_655, // sfix19_En18 
  input [18:0] Wgt_5_656, // sfix19_En18 
  input [18:0] Wgt_5_657, // sfix19_En18 
  input [18:0] Wgt_5_658, // sfix19_En18 
  input [18:0] Wgt_5_659, // sfix19_En18 
  input [18:0] Wgt_5_660, // sfix19_En18 
  input [18:0] Wgt_5_661, // sfix19_En18 
  input [18:0] Wgt_5_662, // sfix19_En18 
  input [18:0] Wgt_5_663, // sfix19_En18 
  input [18:0] Wgt_5_664, // sfix19_En18 
  input [18:0] Wgt_5_665, // sfix19_En18 
  input [18:0] Wgt_5_666, // sfix19_En18 
  input [18:0] Wgt_5_667, // sfix19_En18 
  input [18:0] Wgt_5_668, // sfix19_En18 
  input [18:0] Wgt_5_669, // sfix19_En18 
  input [18:0] Wgt_5_670, // sfix19_En18 
  input [18:0] Wgt_5_671, // sfix19_En18 
  input [18:0] Wgt_5_672, // sfix19_En18 
  input [18:0] Wgt_5_673, // sfix19_En18 
  input [18:0] Wgt_5_674, // sfix19_En18 
  input [18:0] Wgt_5_675, // sfix19_En18 
  input [18:0] Wgt_5_676, // sfix19_En18 
  input [18:0] Wgt_5_677, // sfix19_En18 
  input [18:0] Wgt_5_678, // sfix19_En18 
  input [18:0] Wgt_5_679, // sfix19_En18 
  input [18:0] Wgt_5_680, // sfix19_En18 
  input [18:0] Wgt_5_681, // sfix19_En18 
  input [18:0] Wgt_5_682, // sfix19_En18 
  input [18:0] Wgt_5_683, // sfix19_En18 
  input [18:0] Wgt_5_684, // sfix19_En18 
  input [18:0] Wgt_5_685, // sfix19_En18 
  input [18:0] Wgt_5_686, // sfix19_En18 
  input [18:0] Wgt_5_687, // sfix19_En18 
  input [18:0] Wgt_5_688, // sfix19_En18 
  input [18:0] Wgt_5_689, // sfix19_En18 
  input [18:0] Wgt_5_690, // sfix19_En18 
  input [18:0] Wgt_5_691, // sfix19_En18 
  input [18:0] Wgt_5_692, // sfix19_En18 
  input [18:0] Wgt_5_693, // sfix19_En18 
  input [18:0] Wgt_5_694, // sfix19_En18 
  input [18:0] Wgt_5_695, // sfix19_En18 
  input [18:0] Wgt_5_696, // sfix19_En18 
  input [18:0] Wgt_5_697, // sfix19_En18 
  input [18:0] Wgt_5_698, // sfix19_En18 
  input [18:0] Wgt_5_699, // sfix19_En18 
  input [18:0] Wgt_5_700, // sfix19_En18 
  input [18:0] Wgt_5_701, // sfix19_En18 
  input [18:0] Wgt_5_702, // sfix19_En18 
  input [18:0] Wgt_5_703, // sfix19_En18 
  input [18:0] Wgt_5_704, // sfix19_En18 
  input [18:0] Wgt_5_705, // sfix19_En18 
  input [18:0] Wgt_5_706, // sfix19_En18 
  input [18:0] Wgt_5_707, // sfix19_En18 
  input [18:0] Wgt_5_708, // sfix19_En18 
  input [18:0] Wgt_5_709, // sfix19_En18 
  input [18:0] Wgt_5_710, // sfix19_En18 
  input [18:0] Wgt_5_711, // sfix19_En18 
  input [18:0] Wgt_5_712, // sfix19_En18 
  input [18:0] Wgt_5_713, // sfix19_En18 
  input [18:0] Wgt_5_714, // sfix19_En18 
  input [18:0] Wgt_5_715, // sfix19_En18 
  input [18:0] Wgt_5_716, // sfix19_En18 
  input [18:0] Wgt_5_717, // sfix19_En18 
  input [18:0] Wgt_5_718, // sfix19_En18 
  input [18:0] Wgt_5_719, // sfix19_En18 
  input [18:0] Wgt_5_720, // sfix19_En18 
  input [18:0] Wgt_5_721, // sfix19_En18 
  input [18:0] Wgt_5_722, // sfix19_En18 
  input [18:0] Wgt_5_723, // sfix19_En18 
  input [18:0] Wgt_5_724, // sfix19_En18 
  input [18:0] Wgt_5_725, // sfix19_En18 
  input [18:0] Wgt_5_726, // sfix19_En18 
  input [18:0] Wgt_5_727, // sfix19_En18 
  input [18:0] Wgt_5_728, // sfix19_En18 
  input [18:0] Wgt_5_729, // sfix19_En18 
  input [18:0] Wgt_5_730, // sfix19_En18 
  input [18:0] Wgt_5_731, // sfix19_En18 
  input [18:0] Wgt_5_732, // sfix19_En18 
  input [18:0] Wgt_5_733, // sfix19_En18 
  input [18:0] Wgt_5_734, // sfix19_En18 
  input [18:0] Wgt_5_735, // sfix19_En18 
  input [18:0] Wgt_5_736, // sfix19_En18 
  input [18:0] Wgt_5_737, // sfix19_En18 
  input [18:0] Wgt_5_738, // sfix19_En18 
  input [18:0] Wgt_5_739, // sfix19_En18 
  input [18:0] Wgt_5_740, // sfix19_En18 
  input [18:0] Wgt_5_741, // sfix19_En18 
  input [18:0] Wgt_5_742, // sfix19_En18 
  input [18:0] Wgt_5_743, // sfix19_En18 
  input [18:0] Wgt_5_744, // sfix19_En18 
  input [18:0] Wgt_5_745, // sfix19_En18 
  input [18:0] Wgt_5_746, // sfix19_En18 
  input [18:0] Wgt_5_747, // sfix19_En18 
  input [18:0] Wgt_5_748, // sfix19_En18 
  input [18:0] Wgt_5_749, // sfix19_En18 
  input [18:0] Wgt_5_750, // sfix19_En18 
  input [18:0] Wgt_5_751, // sfix19_En18 
  input [18:0] Wgt_5_752, // sfix19_En18 
  input [18:0] Wgt_5_753, // sfix19_En18 
  input [18:0] Wgt_5_754, // sfix19_En18 
  input [18:0] Wgt_5_755, // sfix19_En18 
  input [18:0] Wgt_5_756, // sfix19_En18 
  input [18:0] Wgt_5_757, // sfix19_En18 
  input [18:0] Wgt_5_758, // sfix19_En18 
  input [18:0] Wgt_5_759, // sfix19_En18 
  input [18:0] Wgt_5_760, // sfix19_En18 
  input [18:0] Wgt_5_761, // sfix19_En18 
  input [18:0] Wgt_5_762, // sfix19_En18 
  input [18:0] Wgt_5_763, // sfix19_En18 
  input [18:0] Wgt_5_764, // sfix19_En18 
  input [18:0] Wgt_5_765, // sfix19_En18 
  input [18:0] Wgt_5_766, // sfix19_En18 
  input [18:0] Wgt_5_767, // sfix19_En18 
  input [18:0] Wgt_5_768, // sfix19_En18 
  input [18:0] Wgt_5_769, // sfix19_En18 
  input [18:0] Wgt_5_770, // sfix19_En18 
  input [18:0] Wgt_5_771, // sfix19_En18 
  input [18:0] Wgt_5_772, // sfix19_En18 
  input [18:0] Wgt_5_773, // sfix19_En18 
  input [18:0] Wgt_5_774, // sfix19_En18 
  input [18:0] Wgt_5_775, // sfix19_En18 
  input [18:0] Wgt_5_776, // sfix19_En18 
  input [18:0] Wgt_5_777, // sfix19_En18 
  input [18:0] Wgt_5_778, // sfix19_En18 
  input [18:0] Wgt_5_779, // sfix19_En18 
  input [18:0] Wgt_5_780, // sfix19_En18 
  input [18:0] Wgt_5_781, // sfix19_En18 
  input [18:0] Wgt_5_782, // sfix19_En18 
  input [18:0] Wgt_5_783, // sfix19_En18 
  input [18:0] Wgt_5_784, // sfix19_En18 
  input [18:0] Wgt_6_0, // sfix19_En18 
  input [18:0] Wgt_6_1, // sfix19_En18 
  input [18:0] Wgt_6_2, // sfix19_En18 
  input [18:0] Wgt_6_3, // sfix19_En18 
  input [18:0] Wgt_6_4, // sfix19_En18 
  input [18:0] Wgt_6_5, // sfix19_En18 
  input [18:0] Wgt_6_6, // sfix19_En18 
  input [18:0] Wgt_6_7, // sfix19_En18 
  input [18:0] Wgt_6_8, // sfix19_En18 
  input [18:0] Wgt_6_9, // sfix19_En18 
  input [18:0] Wgt_6_10, // sfix19_En18 
  input [18:0] Wgt_6_11, // sfix19_En18 
  input [18:0] Wgt_6_12, // sfix19_En18 
  input [18:0] Wgt_6_13, // sfix19_En18 
  input [18:0] Wgt_6_14, // sfix19_En18 
  input [18:0] Wgt_6_15, // sfix19_En18 
  input [18:0] Wgt_6_16, // sfix19_En18 
  input [18:0] Wgt_6_17, // sfix19_En18 
  input [18:0] Wgt_6_18, // sfix19_En18 
  input [18:0] Wgt_6_19, // sfix19_En18 
  input [18:0] Wgt_6_20, // sfix19_En18 
  input [18:0] Wgt_6_21, // sfix19_En18 
  input [18:0] Wgt_6_22, // sfix19_En18 
  input [18:0] Wgt_6_23, // sfix19_En18 
  input [18:0] Wgt_6_24, // sfix19_En18 
  input [18:0] Wgt_6_25, // sfix19_En18 
  input [18:0] Wgt_6_26, // sfix19_En18 
  input [18:0] Wgt_6_27, // sfix19_En18 
  input [18:0] Wgt_6_28, // sfix19_En18 
  input [18:0] Wgt_6_29, // sfix19_En18 
  input [18:0] Wgt_6_30, // sfix19_En18 
  input [18:0] Wgt_6_31, // sfix19_En18 
  input [18:0] Wgt_6_32, // sfix19_En18 
  input [18:0] Wgt_6_33, // sfix19_En18 
  input [18:0] Wgt_6_34, // sfix19_En18 
  input [18:0] Wgt_6_35, // sfix19_En18 
  input [18:0] Wgt_6_36, // sfix19_En18 
  input [18:0] Wgt_6_37, // sfix19_En18 
  input [18:0] Wgt_6_38, // sfix19_En18 
  input [18:0] Wgt_6_39, // sfix19_En18 
  input [18:0] Wgt_6_40, // sfix19_En18 
  input [18:0] Wgt_6_41, // sfix19_En18 
  input [18:0] Wgt_6_42, // sfix19_En18 
  input [18:0] Wgt_6_43, // sfix19_En18 
  input [18:0] Wgt_6_44, // sfix19_En18 
  input [18:0] Wgt_6_45, // sfix19_En18 
  input [18:0] Wgt_6_46, // sfix19_En18 
  input [18:0] Wgt_6_47, // sfix19_En18 
  input [18:0] Wgt_6_48, // sfix19_En18 
  input [18:0] Wgt_6_49, // sfix19_En18 
  input [18:0] Wgt_6_50, // sfix19_En18 
  input [18:0] Wgt_6_51, // sfix19_En18 
  input [18:0] Wgt_6_52, // sfix19_En18 
  input [18:0] Wgt_6_53, // sfix19_En18 
  input [18:0] Wgt_6_54, // sfix19_En18 
  input [18:0] Wgt_6_55, // sfix19_En18 
  input [18:0] Wgt_6_56, // sfix19_En18 
  input [18:0] Wgt_6_57, // sfix19_En18 
  input [18:0] Wgt_6_58, // sfix19_En18 
  input [18:0] Wgt_6_59, // sfix19_En18 
  input [18:0] Wgt_6_60, // sfix19_En18 
  input [18:0] Wgt_6_61, // sfix19_En18 
  input [18:0] Wgt_6_62, // sfix19_En18 
  input [18:0] Wgt_6_63, // sfix19_En18 
  input [18:0] Wgt_6_64, // sfix19_En18 
  input [18:0] Wgt_6_65, // sfix19_En18 
  input [18:0] Wgt_6_66, // sfix19_En18 
  input [18:0] Wgt_6_67, // sfix19_En18 
  input [18:0] Wgt_6_68, // sfix19_En18 
  input [18:0] Wgt_6_69, // sfix19_En18 
  input [18:0] Wgt_6_70, // sfix19_En18 
  input [18:0] Wgt_6_71, // sfix19_En18 
  input [18:0] Wgt_6_72, // sfix19_En18 
  input [18:0] Wgt_6_73, // sfix19_En18 
  input [18:0] Wgt_6_74, // sfix19_En18 
  input [18:0] Wgt_6_75, // sfix19_En18 
  input [18:0] Wgt_6_76, // sfix19_En18 
  input [18:0] Wgt_6_77, // sfix19_En18 
  input [18:0] Wgt_6_78, // sfix19_En18 
  input [18:0] Wgt_6_79, // sfix19_En18 
  input [18:0] Wgt_6_80, // sfix19_En18 
  input [18:0] Wgt_6_81, // sfix19_En18 
  input [18:0] Wgt_6_82, // sfix19_En18 
  input [18:0] Wgt_6_83, // sfix19_En18 
  input [18:0] Wgt_6_84, // sfix19_En18 
  input [18:0] Wgt_6_85, // sfix19_En18 
  input [18:0] Wgt_6_86, // sfix19_En18 
  input [18:0] Wgt_6_87, // sfix19_En18 
  input [18:0] Wgt_6_88, // sfix19_En18 
  input [18:0] Wgt_6_89, // sfix19_En18 
  input [18:0] Wgt_6_90, // sfix19_En18 
  input [18:0] Wgt_6_91, // sfix19_En18 
  input [18:0] Wgt_6_92, // sfix19_En18 
  input [18:0] Wgt_6_93, // sfix19_En18 
  input [18:0] Wgt_6_94, // sfix19_En18 
  input [18:0] Wgt_6_95, // sfix19_En18 
  input [18:0] Wgt_6_96, // sfix19_En18 
  input [18:0] Wgt_6_97, // sfix19_En18 
  input [18:0] Wgt_6_98, // sfix19_En18 
  input [18:0] Wgt_6_99, // sfix19_En18 
  input [18:0] Wgt_6_100, // sfix19_En18 
  input [18:0] Wgt_6_101, // sfix19_En18 
  input [18:0] Wgt_6_102, // sfix19_En18 
  input [18:0] Wgt_6_103, // sfix19_En18 
  input [18:0] Wgt_6_104, // sfix19_En18 
  input [18:0] Wgt_6_105, // sfix19_En18 
  input [18:0] Wgt_6_106, // sfix19_En18 
  input [18:0] Wgt_6_107, // sfix19_En18 
  input [18:0] Wgt_6_108, // sfix19_En18 
  input [18:0] Wgt_6_109, // sfix19_En18 
  input [18:0] Wgt_6_110, // sfix19_En18 
  input [18:0] Wgt_6_111, // sfix19_En18 
  input [18:0] Wgt_6_112, // sfix19_En18 
  input [18:0] Wgt_6_113, // sfix19_En18 
  input [18:0] Wgt_6_114, // sfix19_En18 
  input [18:0] Wgt_6_115, // sfix19_En18 
  input [18:0] Wgt_6_116, // sfix19_En18 
  input [18:0] Wgt_6_117, // sfix19_En18 
  input [18:0] Wgt_6_118, // sfix19_En18 
  input [18:0] Wgt_6_119, // sfix19_En18 
  input [18:0] Wgt_6_120, // sfix19_En18 
  input [18:0] Wgt_6_121, // sfix19_En18 
  input [18:0] Wgt_6_122, // sfix19_En18 
  input [18:0] Wgt_6_123, // sfix19_En18 
  input [18:0] Wgt_6_124, // sfix19_En18 
  input [18:0] Wgt_6_125, // sfix19_En18 
  input [18:0] Wgt_6_126, // sfix19_En18 
  input [18:0] Wgt_6_127, // sfix19_En18 
  input [18:0] Wgt_6_128, // sfix19_En18 
  input [18:0] Wgt_6_129, // sfix19_En18 
  input [18:0] Wgt_6_130, // sfix19_En18 
  input [18:0] Wgt_6_131, // sfix19_En18 
  input [18:0] Wgt_6_132, // sfix19_En18 
  input [18:0] Wgt_6_133, // sfix19_En18 
  input [18:0] Wgt_6_134, // sfix19_En18 
  input [18:0] Wgt_6_135, // sfix19_En18 
  input [18:0] Wgt_6_136, // sfix19_En18 
  input [18:0] Wgt_6_137, // sfix19_En18 
  input [18:0] Wgt_6_138, // sfix19_En18 
  input [18:0] Wgt_6_139, // sfix19_En18 
  input [18:0] Wgt_6_140, // sfix19_En18 
  input [18:0] Wgt_6_141, // sfix19_En18 
  input [18:0] Wgt_6_142, // sfix19_En18 
  input [18:0] Wgt_6_143, // sfix19_En18 
  input [18:0] Wgt_6_144, // sfix19_En18 
  input [18:0] Wgt_6_145, // sfix19_En18 
  input [18:0] Wgt_6_146, // sfix19_En18 
  input [18:0] Wgt_6_147, // sfix19_En18 
  input [18:0] Wgt_6_148, // sfix19_En18 
  input [18:0] Wgt_6_149, // sfix19_En18 
  input [18:0] Wgt_6_150, // sfix19_En18 
  input [18:0] Wgt_6_151, // sfix19_En18 
  input [18:0] Wgt_6_152, // sfix19_En18 
  input [18:0] Wgt_6_153, // sfix19_En18 
  input [18:0] Wgt_6_154, // sfix19_En18 
  input [18:0] Wgt_6_155, // sfix19_En18 
  input [18:0] Wgt_6_156, // sfix19_En18 
  input [18:0] Wgt_6_157, // sfix19_En18 
  input [18:0] Wgt_6_158, // sfix19_En18 
  input [18:0] Wgt_6_159, // sfix19_En18 
  input [18:0] Wgt_6_160, // sfix19_En18 
  input [18:0] Wgt_6_161, // sfix19_En18 
  input [18:0] Wgt_6_162, // sfix19_En18 
  input [18:0] Wgt_6_163, // sfix19_En18 
  input [18:0] Wgt_6_164, // sfix19_En18 
  input [18:0] Wgt_6_165, // sfix19_En18 
  input [18:0] Wgt_6_166, // sfix19_En18 
  input [18:0] Wgt_6_167, // sfix19_En18 
  input [18:0] Wgt_6_168, // sfix19_En18 
  input [18:0] Wgt_6_169, // sfix19_En18 
  input [18:0] Wgt_6_170, // sfix19_En18 
  input [18:0] Wgt_6_171, // sfix19_En18 
  input [18:0] Wgt_6_172, // sfix19_En18 
  input [18:0] Wgt_6_173, // sfix19_En18 
  input [18:0] Wgt_6_174, // sfix19_En18 
  input [18:0] Wgt_6_175, // sfix19_En18 
  input [18:0] Wgt_6_176, // sfix19_En18 
  input [18:0] Wgt_6_177, // sfix19_En18 
  input [18:0] Wgt_6_178, // sfix19_En18 
  input [18:0] Wgt_6_179, // sfix19_En18 
  input [18:0] Wgt_6_180, // sfix19_En18 
  input [18:0] Wgt_6_181, // sfix19_En18 
  input [18:0] Wgt_6_182, // sfix19_En18 
  input [18:0] Wgt_6_183, // sfix19_En18 
  input [18:0] Wgt_6_184, // sfix19_En18 
  input [18:0] Wgt_6_185, // sfix19_En18 
  input [18:0] Wgt_6_186, // sfix19_En18 
  input [18:0] Wgt_6_187, // sfix19_En18 
  input [18:0] Wgt_6_188, // sfix19_En18 
  input [18:0] Wgt_6_189, // sfix19_En18 
  input [18:0] Wgt_6_190, // sfix19_En18 
  input [18:0] Wgt_6_191, // sfix19_En18 
  input [18:0] Wgt_6_192, // sfix19_En18 
  input [18:0] Wgt_6_193, // sfix19_En18 
  input [18:0] Wgt_6_194, // sfix19_En18 
  input [18:0] Wgt_6_195, // sfix19_En18 
  input [18:0] Wgt_6_196, // sfix19_En18 
  input [18:0] Wgt_6_197, // sfix19_En18 
  input [18:0] Wgt_6_198, // sfix19_En18 
  input [18:0] Wgt_6_199, // sfix19_En18 
  input [18:0] Wgt_6_200, // sfix19_En18 
  input [18:0] Wgt_6_201, // sfix19_En18 
  input [18:0] Wgt_6_202, // sfix19_En18 
  input [18:0] Wgt_6_203, // sfix19_En18 
  input [18:0] Wgt_6_204, // sfix19_En18 
  input [18:0] Wgt_6_205, // sfix19_En18 
  input [18:0] Wgt_6_206, // sfix19_En18 
  input [18:0] Wgt_6_207, // sfix19_En18 
  input [18:0] Wgt_6_208, // sfix19_En18 
  input [18:0] Wgt_6_209, // sfix19_En18 
  input [18:0] Wgt_6_210, // sfix19_En18 
  input [18:0] Wgt_6_211, // sfix19_En18 
  input [18:0] Wgt_6_212, // sfix19_En18 
  input [18:0] Wgt_6_213, // sfix19_En18 
  input [18:0] Wgt_6_214, // sfix19_En18 
  input [18:0] Wgt_6_215, // sfix19_En18 
  input [18:0] Wgt_6_216, // sfix19_En18 
  input [18:0] Wgt_6_217, // sfix19_En18 
  input [18:0] Wgt_6_218, // sfix19_En18 
  input [18:0] Wgt_6_219, // sfix19_En18 
  input [18:0] Wgt_6_220, // sfix19_En18 
  input [18:0] Wgt_6_221, // sfix19_En18 
  input [18:0] Wgt_6_222, // sfix19_En18 
  input [18:0] Wgt_6_223, // sfix19_En18 
  input [18:0] Wgt_6_224, // sfix19_En18 
  input [18:0] Wgt_6_225, // sfix19_En18 
  input [18:0] Wgt_6_226, // sfix19_En18 
  input [18:0] Wgt_6_227, // sfix19_En18 
  input [18:0] Wgt_6_228, // sfix19_En18 
  input [18:0] Wgt_6_229, // sfix19_En18 
  input [18:0] Wgt_6_230, // sfix19_En18 
  input [18:0] Wgt_6_231, // sfix19_En18 
  input [18:0] Wgt_6_232, // sfix19_En18 
  input [18:0] Wgt_6_233, // sfix19_En18 
  input [18:0] Wgt_6_234, // sfix19_En18 
  input [18:0] Wgt_6_235, // sfix19_En18 
  input [18:0] Wgt_6_236, // sfix19_En18 
  input [18:0] Wgt_6_237, // sfix19_En18 
  input [18:0] Wgt_6_238, // sfix19_En18 
  input [18:0] Wgt_6_239, // sfix19_En18 
  input [18:0] Wgt_6_240, // sfix19_En18 
  input [18:0] Wgt_6_241, // sfix19_En18 
  input [18:0] Wgt_6_242, // sfix19_En18 
  input [18:0] Wgt_6_243, // sfix19_En18 
  input [18:0] Wgt_6_244, // sfix19_En18 
  input [18:0] Wgt_6_245, // sfix19_En18 
  input [18:0] Wgt_6_246, // sfix19_En18 
  input [18:0] Wgt_6_247, // sfix19_En18 
  input [18:0] Wgt_6_248, // sfix19_En18 
  input [18:0] Wgt_6_249, // sfix19_En18 
  input [18:0] Wgt_6_250, // sfix19_En18 
  input [18:0] Wgt_6_251, // sfix19_En18 
  input [18:0] Wgt_6_252, // sfix19_En18 
  input [18:0] Wgt_6_253, // sfix19_En18 
  input [18:0] Wgt_6_254, // sfix19_En18 
  input [18:0] Wgt_6_255, // sfix19_En18 
  input [18:0] Wgt_6_256, // sfix19_En18 
  input [18:0] Wgt_6_257, // sfix19_En18 
  input [18:0] Wgt_6_258, // sfix19_En18 
  input [18:0] Wgt_6_259, // sfix19_En18 
  input [18:0] Wgt_6_260, // sfix19_En18 
  input [18:0] Wgt_6_261, // sfix19_En18 
  input [18:0] Wgt_6_262, // sfix19_En18 
  input [18:0] Wgt_6_263, // sfix19_En18 
  input [18:0] Wgt_6_264, // sfix19_En18 
  input [18:0] Wgt_6_265, // sfix19_En18 
  input [18:0] Wgt_6_266, // sfix19_En18 
  input [18:0] Wgt_6_267, // sfix19_En18 
  input [18:0] Wgt_6_268, // sfix19_En18 
  input [18:0] Wgt_6_269, // sfix19_En18 
  input [18:0] Wgt_6_270, // sfix19_En18 
  input [18:0] Wgt_6_271, // sfix19_En18 
  input [18:0] Wgt_6_272, // sfix19_En18 
  input [18:0] Wgt_6_273, // sfix19_En18 
  input [18:0] Wgt_6_274, // sfix19_En18 
  input [18:0] Wgt_6_275, // sfix19_En18 
  input [18:0] Wgt_6_276, // sfix19_En18 
  input [18:0] Wgt_6_277, // sfix19_En18 
  input [18:0] Wgt_6_278, // sfix19_En18 
  input [18:0] Wgt_6_279, // sfix19_En18 
  input [18:0] Wgt_6_280, // sfix19_En18 
  input [18:0] Wgt_6_281, // sfix19_En18 
  input [18:0] Wgt_6_282, // sfix19_En18 
  input [18:0] Wgt_6_283, // sfix19_En18 
  input [18:0] Wgt_6_284, // sfix19_En18 
  input [18:0] Wgt_6_285, // sfix19_En18 
  input [18:0] Wgt_6_286, // sfix19_En18 
  input [18:0] Wgt_6_287, // sfix19_En18 
  input [18:0] Wgt_6_288, // sfix19_En18 
  input [18:0] Wgt_6_289, // sfix19_En18 
  input [18:0] Wgt_6_290, // sfix19_En18 
  input [18:0] Wgt_6_291, // sfix19_En18 
  input [18:0] Wgt_6_292, // sfix19_En18 
  input [18:0] Wgt_6_293, // sfix19_En18 
  input [18:0] Wgt_6_294, // sfix19_En18 
  input [18:0] Wgt_6_295, // sfix19_En18 
  input [18:0] Wgt_6_296, // sfix19_En18 
  input [18:0] Wgt_6_297, // sfix19_En18 
  input [18:0] Wgt_6_298, // sfix19_En18 
  input [18:0] Wgt_6_299, // sfix19_En18 
  input [18:0] Wgt_6_300, // sfix19_En18 
  input [18:0] Wgt_6_301, // sfix19_En18 
  input [18:0] Wgt_6_302, // sfix19_En18 
  input [18:0] Wgt_6_303, // sfix19_En18 
  input [18:0] Wgt_6_304, // sfix19_En18 
  input [18:0] Wgt_6_305, // sfix19_En18 
  input [18:0] Wgt_6_306, // sfix19_En18 
  input [18:0] Wgt_6_307, // sfix19_En18 
  input [18:0] Wgt_6_308, // sfix19_En18 
  input [18:0] Wgt_6_309, // sfix19_En18 
  input [18:0] Wgt_6_310, // sfix19_En18 
  input [18:0] Wgt_6_311, // sfix19_En18 
  input [18:0] Wgt_6_312, // sfix19_En18 
  input [18:0] Wgt_6_313, // sfix19_En18 
  input [18:0] Wgt_6_314, // sfix19_En18 
  input [18:0] Wgt_6_315, // sfix19_En18 
  input [18:0] Wgt_6_316, // sfix19_En18 
  input [18:0] Wgt_6_317, // sfix19_En18 
  input [18:0] Wgt_6_318, // sfix19_En18 
  input [18:0] Wgt_6_319, // sfix19_En18 
  input [18:0] Wgt_6_320, // sfix19_En18 
  input [18:0] Wgt_6_321, // sfix19_En18 
  input [18:0] Wgt_6_322, // sfix19_En18 
  input [18:0] Wgt_6_323, // sfix19_En18 
  input [18:0] Wgt_6_324, // sfix19_En18 
  input [18:0] Wgt_6_325, // sfix19_En18 
  input [18:0] Wgt_6_326, // sfix19_En18 
  input [18:0] Wgt_6_327, // sfix19_En18 
  input [18:0] Wgt_6_328, // sfix19_En18 
  input [18:0] Wgt_6_329, // sfix19_En18 
  input [18:0] Wgt_6_330, // sfix19_En18 
  input [18:0] Wgt_6_331, // sfix19_En18 
  input [18:0] Wgt_6_332, // sfix19_En18 
  input [18:0] Wgt_6_333, // sfix19_En18 
  input [18:0] Wgt_6_334, // sfix19_En18 
  input [18:0] Wgt_6_335, // sfix19_En18 
  input [18:0] Wgt_6_336, // sfix19_En18 
  input [18:0] Wgt_6_337, // sfix19_En18 
  input [18:0] Wgt_6_338, // sfix19_En18 
  input [18:0] Wgt_6_339, // sfix19_En18 
  input [18:0] Wgt_6_340, // sfix19_En18 
  input [18:0] Wgt_6_341, // sfix19_En18 
  input [18:0] Wgt_6_342, // sfix19_En18 
  input [18:0] Wgt_6_343, // sfix19_En18 
  input [18:0] Wgt_6_344, // sfix19_En18 
  input [18:0] Wgt_6_345, // sfix19_En18 
  input [18:0] Wgt_6_346, // sfix19_En18 
  input [18:0] Wgt_6_347, // sfix19_En18 
  input [18:0] Wgt_6_348, // sfix19_En18 
  input [18:0] Wgt_6_349, // sfix19_En18 
  input [18:0] Wgt_6_350, // sfix19_En18 
  input [18:0] Wgt_6_351, // sfix19_En18 
  input [18:0] Wgt_6_352, // sfix19_En18 
  input [18:0] Wgt_6_353, // sfix19_En18 
  input [18:0] Wgt_6_354, // sfix19_En18 
  input [18:0] Wgt_6_355, // sfix19_En18 
  input [18:0] Wgt_6_356, // sfix19_En18 
  input [18:0] Wgt_6_357, // sfix19_En18 
  input [18:0] Wgt_6_358, // sfix19_En18 
  input [18:0] Wgt_6_359, // sfix19_En18 
  input [18:0] Wgt_6_360, // sfix19_En18 
  input [18:0] Wgt_6_361, // sfix19_En18 
  input [18:0] Wgt_6_362, // sfix19_En18 
  input [18:0] Wgt_6_363, // sfix19_En18 
  input [18:0] Wgt_6_364, // sfix19_En18 
  input [18:0] Wgt_6_365, // sfix19_En18 
  input [18:0] Wgt_6_366, // sfix19_En18 
  input [18:0] Wgt_6_367, // sfix19_En18 
  input [18:0] Wgt_6_368, // sfix19_En18 
  input [18:0] Wgt_6_369, // sfix19_En18 
  input [18:0] Wgt_6_370, // sfix19_En18 
  input [18:0] Wgt_6_371, // sfix19_En18 
  input [18:0] Wgt_6_372, // sfix19_En18 
  input [18:0] Wgt_6_373, // sfix19_En18 
  input [18:0] Wgt_6_374, // sfix19_En18 
  input [18:0] Wgt_6_375, // sfix19_En18 
  input [18:0] Wgt_6_376, // sfix19_En18 
  input [18:0] Wgt_6_377, // sfix19_En18 
  input [18:0] Wgt_6_378, // sfix19_En18 
  input [18:0] Wgt_6_379, // sfix19_En18 
  input [18:0] Wgt_6_380, // sfix19_En18 
  input [18:0] Wgt_6_381, // sfix19_En18 
  input [18:0] Wgt_6_382, // sfix19_En18 
  input [18:0] Wgt_6_383, // sfix19_En18 
  input [18:0] Wgt_6_384, // sfix19_En18 
  input [18:0] Wgt_6_385, // sfix19_En18 
  input [18:0] Wgt_6_386, // sfix19_En18 
  input [18:0] Wgt_6_387, // sfix19_En18 
  input [18:0] Wgt_6_388, // sfix19_En18 
  input [18:0] Wgt_6_389, // sfix19_En18 
  input [18:0] Wgt_6_390, // sfix19_En18 
  input [18:0] Wgt_6_391, // sfix19_En18 
  input [18:0] Wgt_6_392, // sfix19_En18 
  input [18:0] Wgt_6_393, // sfix19_En18 
  input [18:0] Wgt_6_394, // sfix19_En18 
  input [18:0] Wgt_6_395, // sfix19_En18 
  input [18:0] Wgt_6_396, // sfix19_En18 
  input [18:0] Wgt_6_397, // sfix19_En18 
  input [18:0] Wgt_6_398, // sfix19_En18 
  input [18:0] Wgt_6_399, // sfix19_En18 
  input [18:0] Wgt_6_400, // sfix19_En18 
  input [18:0] Wgt_6_401, // sfix19_En18 
  input [18:0] Wgt_6_402, // sfix19_En18 
  input [18:0] Wgt_6_403, // sfix19_En18 
  input [18:0] Wgt_6_404, // sfix19_En18 
  input [18:0] Wgt_6_405, // sfix19_En18 
  input [18:0] Wgt_6_406, // sfix19_En18 
  input [18:0] Wgt_6_407, // sfix19_En18 
  input [18:0] Wgt_6_408, // sfix19_En18 
  input [18:0] Wgt_6_409, // sfix19_En18 
  input [18:0] Wgt_6_410, // sfix19_En18 
  input [18:0] Wgt_6_411, // sfix19_En18 
  input [18:0] Wgt_6_412, // sfix19_En18 
  input [18:0] Wgt_6_413, // sfix19_En18 
  input [18:0] Wgt_6_414, // sfix19_En18 
  input [18:0] Wgt_6_415, // sfix19_En18 
  input [18:0] Wgt_6_416, // sfix19_En18 
  input [18:0] Wgt_6_417, // sfix19_En18 
  input [18:0] Wgt_6_418, // sfix19_En18 
  input [18:0] Wgt_6_419, // sfix19_En18 
  input [18:0] Wgt_6_420, // sfix19_En18 
  input [18:0] Wgt_6_421, // sfix19_En18 
  input [18:0] Wgt_6_422, // sfix19_En18 
  input [18:0] Wgt_6_423, // sfix19_En18 
  input [18:0] Wgt_6_424, // sfix19_En18 
  input [18:0] Wgt_6_425, // sfix19_En18 
  input [18:0] Wgt_6_426, // sfix19_En18 
  input [18:0] Wgt_6_427, // sfix19_En18 
  input [18:0] Wgt_6_428, // sfix19_En18 
  input [18:0] Wgt_6_429, // sfix19_En18 
  input [18:0] Wgt_6_430, // sfix19_En18 
  input [18:0] Wgt_6_431, // sfix19_En18 
  input [18:0] Wgt_6_432, // sfix19_En18 
  input [18:0] Wgt_6_433, // sfix19_En18 
  input [18:0] Wgt_6_434, // sfix19_En18 
  input [18:0] Wgt_6_435, // sfix19_En18 
  input [18:0] Wgt_6_436, // sfix19_En18 
  input [18:0] Wgt_6_437, // sfix19_En18 
  input [18:0] Wgt_6_438, // sfix19_En18 
  input [18:0] Wgt_6_439, // sfix19_En18 
  input [18:0] Wgt_6_440, // sfix19_En18 
  input [18:0] Wgt_6_441, // sfix19_En18 
  input [18:0] Wgt_6_442, // sfix19_En18 
  input [18:0] Wgt_6_443, // sfix19_En18 
  input [18:0] Wgt_6_444, // sfix19_En18 
  input [18:0] Wgt_6_445, // sfix19_En18 
  input [18:0] Wgt_6_446, // sfix19_En18 
  input [18:0] Wgt_6_447, // sfix19_En18 
  input [18:0] Wgt_6_448, // sfix19_En18 
  input [18:0] Wgt_6_449, // sfix19_En18 
  input [18:0] Wgt_6_450, // sfix19_En18 
  input [18:0] Wgt_6_451, // sfix19_En18 
  input [18:0] Wgt_6_452, // sfix19_En18 
  input [18:0] Wgt_6_453, // sfix19_En18 
  input [18:0] Wgt_6_454, // sfix19_En18 
  input [18:0] Wgt_6_455, // sfix19_En18 
  input [18:0] Wgt_6_456, // sfix19_En18 
  input [18:0] Wgt_6_457, // sfix19_En18 
  input [18:0] Wgt_6_458, // sfix19_En18 
  input [18:0] Wgt_6_459, // sfix19_En18 
  input [18:0] Wgt_6_460, // sfix19_En18 
  input [18:0] Wgt_6_461, // sfix19_En18 
  input [18:0] Wgt_6_462, // sfix19_En18 
  input [18:0] Wgt_6_463, // sfix19_En18 
  input [18:0] Wgt_6_464, // sfix19_En18 
  input [18:0] Wgt_6_465, // sfix19_En18 
  input [18:0] Wgt_6_466, // sfix19_En18 
  input [18:0] Wgt_6_467, // sfix19_En18 
  input [18:0] Wgt_6_468, // sfix19_En18 
  input [18:0] Wgt_6_469, // sfix19_En18 
  input [18:0] Wgt_6_470, // sfix19_En18 
  input [18:0] Wgt_6_471, // sfix19_En18 
  input [18:0] Wgt_6_472, // sfix19_En18 
  input [18:0] Wgt_6_473, // sfix19_En18 
  input [18:0] Wgt_6_474, // sfix19_En18 
  input [18:0] Wgt_6_475, // sfix19_En18 
  input [18:0] Wgt_6_476, // sfix19_En18 
  input [18:0] Wgt_6_477, // sfix19_En18 
  input [18:0] Wgt_6_478, // sfix19_En18 
  input [18:0] Wgt_6_479, // sfix19_En18 
  input [18:0] Wgt_6_480, // sfix19_En18 
  input [18:0] Wgt_6_481, // sfix19_En18 
  input [18:0] Wgt_6_482, // sfix19_En18 
  input [18:0] Wgt_6_483, // sfix19_En18 
  input [18:0] Wgt_6_484, // sfix19_En18 
  input [18:0] Wgt_6_485, // sfix19_En18 
  input [18:0] Wgt_6_486, // sfix19_En18 
  input [18:0] Wgt_6_487, // sfix19_En18 
  input [18:0] Wgt_6_488, // sfix19_En18 
  input [18:0] Wgt_6_489, // sfix19_En18 
  input [18:0] Wgt_6_490, // sfix19_En18 
  input [18:0] Wgt_6_491, // sfix19_En18 
  input [18:0] Wgt_6_492, // sfix19_En18 
  input [18:0] Wgt_6_493, // sfix19_En18 
  input [18:0] Wgt_6_494, // sfix19_En18 
  input [18:0] Wgt_6_495, // sfix19_En18 
  input [18:0] Wgt_6_496, // sfix19_En18 
  input [18:0] Wgt_6_497, // sfix19_En18 
  input [18:0] Wgt_6_498, // sfix19_En18 
  input [18:0] Wgt_6_499, // sfix19_En18 
  input [18:0] Wgt_6_500, // sfix19_En18 
  input [18:0] Wgt_6_501, // sfix19_En18 
  input [18:0] Wgt_6_502, // sfix19_En18 
  input [18:0] Wgt_6_503, // sfix19_En18 
  input [18:0] Wgt_6_504, // sfix19_En18 
  input [18:0] Wgt_6_505, // sfix19_En18 
  input [18:0] Wgt_6_506, // sfix19_En18 
  input [18:0] Wgt_6_507, // sfix19_En18 
  input [18:0] Wgt_6_508, // sfix19_En18 
  input [18:0] Wgt_6_509, // sfix19_En18 
  input [18:0] Wgt_6_510, // sfix19_En18 
  input [18:0] Wgt_6_511, // sfix19_En18 
  input [18:0] Wgt_6_512, // sfix19_En18 
  input [18:0] Wgt_6_513, // sfix19_En18 
  input [18:0] Wgt_6_514, // sfix19_En18 
  input [18:0] Wgt_6_515, // sfix19_En18 
  input [18:0] Wgt_6_516, // sfix19_En18 
  input [18:0] Wgt_6_517, // sfix19_En18 
  input [18:0] Wgt_6_518, // sfix19_En18 
  input [18:0] Wgt_6_519, // sfix19_En18 
  input [18:0] Wgt_6_520, // sfix19_En18 
  input [18:0] Wgt_6_521, // sfix19_En18 
  input [18:0] Wgt_6_522, // sfix19_En18 
  input [18:0] Wgt_6_523, // sfix19_En18 
  input [18:0] Wgt_6_524, // sfix19_En18 
  input [18:0] Wgt_6_525, // sfix19_En18 
  input [18:0] Wgt_6_526, // sfix19_En18 
  input [18:0] Wgt_6_527, // sfix19_En18 
  input [18:0] Wgt_6_528, // sfix19_En18 
  input [18:0] Wgt_6_529, // sfix19_En18 
  input [18:0] Wgt_6_530, // sfix19_En18 
  input [18:0] Wgt_6_531, // sfix19_En18 
  input [18:0] Wgt_6_532, // sfix19_En18 
  input [18:0] Wgt_6_533, // sfix19_En18 
  input [18:0] Wgt_6_534, // sfix19_En18 
  input [18:0] Wgt_6_535, // sfix19_En18 
  input [18:0] Wgt_6_536, // sfix19_En18 
  input [18:0] Wgt_6_537, // sfix19_En18 
  input [18:0] Wgt_6_538, // sfix19_En18 
  input [18:0] Wgt_6_539, // sfix19_En18 
  input [18:0] Wgt_6_540, // sfix19_En18 
  input [18:0] Wgt_6_541, // sfix19_En18 
  input [18:0] Wgt_6_542, // sfix19_En18 
  input [18:0] Wgt_6_543, // sfix19_En18 
  input [18:0] Wgt_6_544, // sfix19_En18 
  input [18:0] Wgt_6_545, // sfix19_En18 
  input [18:0] Wgt_6_546, // sfix19_En18 
  input [18:0] Wgt_6_547, // sfix19_En18 
  input [18:0] Wgt_6_548, // sfix19_En18 
  input [18:0] Wgt_6_549, // sfix19_En18 
  input [18:0] Wgt_6_550, // sfix19_En18 
  input [18:0] Wgt_6_551, // sfix19_En18 
  input [18:0] Wgt_6_552, // sfix19_En18 
  input [18:0] Wgt_6_553, // sfix19_En18 
  input [18:0] Wgt_6_554, // sfix19_En18 
  input [18:0] Wgt_6_555, // sfix19_En18 
  input [18:0] Wgt_6_556, // sfix19_En18 
  input [18:0] Wgt_6_557, // sfix19_En18 
  input [18:0] Wgt_6_558, // sfix19_En18 
  input [18:0] Wgt_6_559, // sfix19_En18 
  input [18:0] Wgt_6_560, // sfix19_En18 
  input [18:0] Wgt_6_561, // sfix19_En18 
  input [18:0] Wgt_6_562, // sfix19_En18 
  input [18:0] Wgt_6_563, // sfix19_En18 
  input [18:0] Wgt_6_564, // sfix19_En18 
  input [18:0] Wgt_6_565, // sfix19_En18 
  input [18:0] Wgt_6_566, // sfix19_En18 
  input [18:0] Wgt_6_567, // sfix19_En18 
  input [18:0] Wgt_6_568, // sfix19_En18 
  input [18:0] Wgt_6_569, // sfix19_En18 
  input [18:0] Wgt_6_570, // sfix19_En18 
  input [18:0] Wgt_6_571, // sfix19_En18 
  input [18:0] Wgt_6_572, // sfix19_En18 
  input [18:0] Wgt_6_573, // sfix19_En18 
  input [18:0] Wgt_6_574, // sfix19_En18 
  input [18:0] Wgt_6_575, // sfix19_En18 
  input [18:0] Wgt_6_576, // sfix19_En18 
  input [18:0] Wgt_6_577, // sfix19_En18 
  input [18:0] Wgt_6_578, // sfix19_En18 
  input [18:0] Wgt_6_579, // sfix19_En18 
  input [18:0] Wgt_6_580, // sfix19_En18 
  input [18:0] Wgt_6_581, // sfix19_En18 
  input [18:0] Wgt_6_582, // sfix19_En18 
  input [18:0] Wgt_6_583, // sfix19_En18 
  input [18:0] Wgt_6_584, // sfix19_En18 
  input [18:0] Wgt_6_585, // sfix19_En18 
  input [18:0] Wgt_6_586, // sfix19_En18 
  input [18:0] Wgt_6_587, // sfix19_En18 
  input [18:0] Wgt_6_588, // sfix19_En18 
  input [18:0] Wgt_6_589, // sfix19_En18 
  input [18:0] Wgt_6_590, // sfix19_En18 
  input [18:0] Wgt_6_591, // sfix19_En18 
  input [18:0] Wgt_6_592, // sfix19_En18 
  input [18:0] Wgt_6_593, // sfix19_En18 
  input [18:0] Wgt_6_594, // sfix19_En18 
  input [18:0] Wgt_6_595, // sfix19_En18 
  input [18:0] Wgt_6_596, // sfix19_En18 
  input [18:0] Wgt_6_597, // sfix19_En18 
  input [18:0] Wgt_6_598, // sfix19_En18 
  input [18:0] Wgt_6_599, // sfix19_En18 
  input [18:0] Wgt_6_600, // sfix19_En18 
  input [18:0] Wgt_6_601, // sfix19_En18 
  input [18:0] Wgt_6_602, // sfix19_En18 
  input [18:0] Wgt_6_603, // sfix19_En18 
  input [18:0] Wgt_6_604, // sfix19_En18 
  input [18:0] Wgt_6_605, // sfix19_En18 
  input [18:0] Wgt_6_606, // sfix19_En18 
  input [18:0] Wgt_6_607, // sfix19_En18 
  input [18:0] Wgt_6_608, // sfix19_En18 
  input [18:0] Wgt_6_609, // sfix19_En18 
  input [18:0] Wgt_6_610, // sfix19_En18 
  input [18:0] Wgt_6_611, // sfix19_En18 
  input [18:0] Wgt_6_612, // sfix19_En18 
  input [18:0] Wgt_6_613, // sfix19_En18 
  input [18:0] Wgt_6_614, // sfix19_En18 
  input [18:0] Wgt_6_615, // sfix19_En18 
  input [18:0] Wgt_6_616, // sfix19_En18 
  input [18:0] Wgt_6_617, // sfix19_En18 
  input [18:0] Wgt_6_618, // sfix19_En18 
  input [18:0] Wgt_6_619, // sfix19_En18 
  input [18:0] Wgt_6_620, // sfix19_En18 
  input [18:0] Wgt_6_621, // sfix19_En18 
  input [18:0] Wgt_6_622, // sfix19_En18 
  input [18:0] Wgt_6_623, // sfix19_En18 
  input [18:0] Wgt_6_624, // sfix19_En18 
  input [18:0] Wgt_6_625, // sfix19_En18 
  input [18:0] Wgt_6_626, // sfix19_En18 
  input [18:0] Wgt_6_627, // sfix19_En18 
  input [18:0] Wgt_6_628, // sfix19_En18 
  input [18:0] Wgt_6_629, // sfix19_En18 
  input [18:0] Wgt_6_630, // sfix19_En18 
  input [18:0] Wgt_6_631, // sfix19_En18 
  input [18:0] Wgt_6_632, // sfix19_En18 
  input [18:0] Wgt_6_633, // sfix19_En18 
  input [18:0] Wgt_6_634, // sfix19_En18 
  input [18:0] Wgt_6_635, // sfix19_En18 
  input [18:0] Wgt_6_636, // sfix19_En18 
  input [18:0] Wgt_6_637, // sfix19_En18 
  input [18:0] Wgt_6_638, // sfix19_En18 
  input [18:0] Wgt_6_639, // sfix19_En18 
  input [18:0] Wgt_6_640, // sfix19_En18 
  input [18:0] Wgt_6_641, // sfix19_En18 
  input [18:0] Wgt_6_642, // sfix19_En18 
  input [18:0] Wgt_6_643, // sfix19_En18 
  input [18:0] Wgt_6_644, // sfix19_En18 
  input [18:0] Wgt_6_645, // sfix19_En18 
  input [18:0] Wgt_6_646, // sfix19_En18 
  input [18:0] Wgt_6_647, // sfix19_En18 
  input [18:0] Wgt_6_648, // sfix19_En18 
  input [18:0] Wgt_6_649, // sfix19_En18 
  input [18:0] Wgt_6_650, // sfix19_En18 
  input [18:0] Wgt_6_651, // sfix19_En18 
  input [18:0] Wgt_6_652, // sfix19_En18 
  input [18:0] Wgt_6_653, // sfix19_En18 
  input [18:0] Wgt_6_654, // sfix19_En18 
  input [18:0] Wgt_6_655, // sfix19_En18 
  input [18:0] Wgt_6_656, // sfix19_En18 
  input [18:0] Wgt_6_657, // sfix19_En18 
  input [18:0] Wgt_6_658, // sfix19_En18 
  input [18:0] Wgt_6_659, // sfix19_En18 
  input [18:0] Wgt_6_660, // sfix19_En18 
  input [18:0] Wgt_6_661, // sfix19_En18 
  input [18:0] Wgt_6_662, // sfix19_En18 
  input [18:0] Wgt_6_663, // sfix19_En18 
  input [18:0] Wgt_6_664, // sfix19_En18 
  input [18:0] Wgt_6_665, // sfix19_En18 
  input [18:0] Wgt_6_666, // sfix19_En18 
  input [18:0] Wgt_6_667, // sfix19_En18 
  input [18:0] Wgt_6_668, // sfix19_En18 
  input [18:0] Wgt_6_669, // sfix19_En18 
  input [18:0] Wgt_6_670, // sfix19_En18 
  input [18:0] Wgt_6_671, // sfix19_En18 
  input [18:0] Wgt_6_672, // sfix19_En18 
  input [18:0] Wgt_6_673, // sfix19_En18 
  input [18:0] Wgt_6_674, // sfix19_En18 
  input [18:0] Wgt_6_675, // sfix19_En18 
  input [18:0] Wgt_6_676, // sfix19_En18 
  input [18:0] Wgt_6_677, // sfix19_En18 
  input [18:0] Wgt_6_678, // sfix19_En18 
  input [18:0] Wgt_6_679, // sfix19_En18 
  input [18:0] Wgt_6_680, // sfix19_En18 
  input [18:0] Wgt_6_681, // sfix19_En18 
  input [18:0] Wgt_6_682, // sfix19_En18 
  input [18:0] Wgt_6_683, // sfix19_En18 
  input [18:0] Wgt_6_684, // sfix19_En18 
  input [18:0] Wgt_6_685, // sfix19_En18 
  input [18:0] Wgt_6_686, // sfix19_En18 
  input [18:0] Wgt_6_687, // sfix19_En18 
  input [18:0] Wgt_6_688, // sfix19_En18 
  input [18:0] Wgt_6_689, // sfix19_En18 
  input [18:0] Wgt_6_690, // sfix19_En18 
  input [18:0] Wgt_6_691, // sfix19_En18 
  input [18:0] Wgt_6_692, // sfix19_En18 
  input [18:0] Wgt_6_693, // sfix19_En18 
  input [18:0] Wgt_6_694, // sfix19_En18 
  input [18:0] Wgt_6_695, // sfix19_En18 
  input [18:0] Wgt_6_696, // sfix19_En18 
  input [18:0] Wgt_6_697, // sfix19_En18 
  input [18:0] Wgt_6_698, // sfix19_En18 
  input [18:0] Wgt_6_699, // sfix19_En18 
  input [18:0] Wgt_6_700, // sfix19_En18 
  input [18:0] Wgt_6_701, // sfix19_En18 
  input [18:0] Wgt_6_702, // sfix19_En18 
  input [18:0] Wgt_6_703, // sfix19_En18 
  input [18:0] Wgt_6_704, // sfix19_En18 
  input [18:0] Wgt_6_705, // sfix19_En18 
  input [18:0] Wgt_6_706, // sfix19_En18 
  input [18:0] Wgt_6_707, // sfix19_En18 
  input [18:0] Wgt_6_708, // sfix19_En18 
  input [18:0] Wgt_6_709, // sfix19_En18 
  input [18:0] Wgt_6_710, // sfix19_En18 
  input [18:0] Wgt_6_711, // sfix19_En18 
  input [18:0] Wgt_6_712, // sfix19_En18 
  input [18:0] Wgt_6_713, // sfix19_En18 
  input [18:0] Wgt_6_714, // sfix19_En18 
  input [18:0] Wgt_6_715, // sfix19_En18 
  input [18:0] Wgt_6_716, // sfix19_En18 
  input [18:0] Wgt_6_717, // sfix19_En18 
  input [18:0] Wgt_6_718, // sfix19_En18 
  input [18:0] Wgt_6_719, // sfix19_En18 
  input [18:0] Wgt_6_720, // sfix19_En18 
  input [18:0] Wgt_6_721, // sfix19_En18 
  input [18:0] Wgt_6_722, // sfix19_En18 
  input [18:0] Wgt_6_723, // sfix19_En18 
  input [18:0] Wgt_6_724, // sfix19_En18 
  input [18:0] Wgt_6_725, // sfix19_En18 
  input [18:0] Wgt_6_726, // sfix19_En18 
  input [18:0] Wgt_6_727, // sfix19_En18 
  input [18:0] Wgt_6_728, // sfix19_En18 
  input [18:0] Wgt_6_729, // sfix19_En18 
  input [18:0] Wgt_6_730, // sfix19_En18 
  input [18:0] Wgt_6_731, // sfix19_En18 
  input [18:0] Wgt_6_732, // sfix19_En18 
  input [18:0] Wgt_6_733, // sfix19_En18 
  input [18:0] Wgt_6_734, // sfix19_En18 
  input [18:0] Wgt_6_735, // sfix19_En18 
  input [18:0] Wgt_6_736, // sfix19_En18 
  input [18:0] Wgt_6_737, // sfix19_En18 
  input [18:0] Wgt_6_738, // sfix19_En18 
  input [18:0] Wgt_6_739, // sfix19_En18 
  input [18:0] Wgt_6_740, // sfix19_En18 
  input [18:0] Wgt_6_741, // sfix19_En18 
  input [18:0] Wgt_6_742, // sfix19_En18 
  input [18:0] Wgt_6_743, // sfix19_En18 
  input [18:0] Wgt_6_744, // sfix19_En18 
  input [18:0] Wgt_6_745, // sfix19_En18 
  input [18:0] Wgt_6_746, // sfix19_En18 
  input [18:0] Wgt_6_747, // sfix19_En18 
  input [18:0] Wgt_6_748, // sfix19_En18 
  input [18:0] Wgt_6_749, // sfix19_En18 
  input [18:0] Wgt_6_750, // sfix19_En18 
  input [18:0] Wgt_6_751, // sfix19_En18 
  input [18:0] Wgt_6_752, // sfix19_En18 
  input [18:0] Wgt_6_753, // sfix19_En18 
  input [18:0] Wgt_6_754, // sfix19_En18 
  input [18:0] Wgt_6_755, // sfix19_En18 
  input [18:0] Wgt_6_756, // sfix19_En18 
  input [18:0] Wgt_6_757, // sfix19_En18 
  input [18:0] Wgt_6_758, // sfix19_En18 
  input [18:0] Wgt_6_759, // sfix19_En18 
  input [18:0] Wgt_6_760, // sfix19_En18 
  input [18:0] Wgt_6_761, // sfix19_En18 
  input [18:0] Wgt_6_762, // sfix19_En18 
  input [18:0] Wgt_6_763, // sfix19_En18 
  input [18:0] Wgt_6_764, // sfix19_En18 
  input [18:0] Wgt_6_765, // sfix19_En18 
  input [18:0] Wgt_6_766, // sfix19_En18 
  input [18:0] Wgt_6_767, // sfix19_En18 
  input [18:0] Wgt_6_768, // sfix19_En18 
  input [18:0] Wgt_6_769, // sfix19_En18 
  input [18:0] Wgt_6_770, // sfix19_En18 
  input [18:0] Wgt_6_771, // sfix19_En18 
  input [18:0] Wgt_6_772, // sfix19_En18 
  input [18:0] Wgt_6_773, // sfix19_En18 
  input [18:0] Wgt_6_774, // sfix19_En18 
  input [18:0] Wgt_6_775, // sfix19_En18 
  input [18:0] Wgt_6_776, // sfix19_En18 
  input [18:0] Wgt_6_777, // sfix19_En18 
  input [18:0] Wgt_6_778, // sfix19_En18 
  input [18:0] Wgt_6_779, // sfix19_En18 
  input [18:0] Wgt_6_780, // sfix19_En18 
  input [18:0] Wgt_6_781, // sfix19_En18 
  input [18:0] Wgt_6_782, // sfix19_En18 
  input [18:0] Wgt_6_783, // sfix19_En18 
  input [18:0] Wgt_6_784, // sfix19_En18 
  input [18:0] Wgt_7_0, // sfix19_En18 
  input [18:0] Wgt_7_1, // sfix19_En18 
  input [18:0] Wgt_7_2, // sfix19_En18 
  input [18:0] Wgt_7_3, // sfix19_En18 
  input [18:0] Wgt_7_4, // sfix19_En18 
  input [18:0] Wgt_7_5, // sfix19_En18 
  input [18:0] Wgt_7_6, // sfix19_En18 
  input [18:0] Wgt_7_7, // sfix19_En18 
  input [18:0] Wgt_7_8, // sfix19_En18 
  input [18:0] Wgt_7_9, // sfix19_En18 
  input [18:0] Wgt_7_10, // sfix19_En18 
  input [18:0] Wgt_7_11, // sfix19_En18 
  input [18:0] Wgt_7_12, // sfix19_En18 
  input [18:0] Wgt_7_13, // sfix19_En18 
  input [18:0] Wgt_7_14, // sfix19_En18 
  input [18:0] Wgt_7_15, // sfix19_En18 
  input [18:0] Wgt_7_16, // sfix19_En18 
  input [18:0] Wgt_7_17, // sfix19_En18 
  input [18:0] Wgt_7_18, // sfix19_En18 
  input [18:0] Wgt_7_19, // sfix19_En18 
  input [18:0] Wgt_7_20, // sfix19_En18 
  input [18:0] Wgt_7_21, // sfix19_En18 
  input [18:0] Wgt_7_22, // sfix19_En18 
  input [18:0] Wgt_7_23, // sfix19_En18 
  input [18:0] Wgt_7_24, // sfix19_En18 
  input [18:0] Wgt_7_25, // sfix19_En18 
  input [18:0] Wgt_7_26, // sfix19_En18 
  input [18:0] Wgt_7_27, // sfix19_En18 
  input [18:0] Wgt_7_28, // sfix19_En18 
  input [18:0] Wgt_7_29, // sfix19_En18 
  input [18:0] Wgt_7_30, // sfix19_En18 
  input [18:0] Wgt_7_31, // sfix19_En18 
  input [18:0] Wgt_7_32, // sfix19_En18 
  input [18:0] Wgt_7_33, // sfix19_En18 
  input [18:0] Wgt_7_34, // sfix19_En18 
  input [18:0] Wgt_7_35, // sfix19_En18 
  input [18:0] Wgt_7_36, // sfix19_En18 
  input [18:0] Wgt_7_37, // sfix19_En18 
  input [18:0] Wgt_7_38, // sfix19_En18 
  input [18:0] Wgt_7_39, // sfix19_En18 
  input [18:0] Wgt_7_40, // sfix19_En18 
  input [18:0] Wgt_7_41, // sfix19_En18 
  input [18:0] Wgt_7_42, // sfix19_En18 
  input [18:0] Wgt_7_43, // sfix19_En18 
  input [18:0] Wgt_7_44, // sfix19_En18 
  input [18:0] Wgt_7_45, // sfix19_En18 
  input [18:0] Wgt_7_46, // sfix19_En18 
  input [18:0] Wgt_7_47, // sfix19_En18 
  input [18:0] Wgt_7_48, // sfix19_En18 
  input [18:0] Wgt_7_49, // sfix19_En18 
  input [18:0] Wgt_7_50, // sfix19_En18 
  input [18:0] Wgt_7_51, // sfix19_En18 
  input [18:0] Wgt_7_52, // sfix19_En18 
  input [18:0] Wgt_7_53, // sfix19_En18 
  input [18:0] Wgt_7_54, // sfix19_En18 
  input [18:0] Wgt_7_55, // sfix19_En18 
  input [18:0] Wgt_7_56, // sfix19_En18 
  input [18:0] Wgt_7_57, // sfix19_En18 
  input [18:0] Wgt_7_58, // sfix19_En18 
  input [18:0] Wgt_7_59, // sfix19_En18 
  input [18:0] Wgt_7_60, // sfix19_En18 
  input [18:0] Wgt_7_61, // sfix19_En18 
  input [18:0] Wgt_7_62, // sfix19_En18 
  input [18:0] Wgt_7_63, // sfix19_En18 
  input [18:0] Wgt_7_64, // sfix19_En18 
  input [18:0] Wgt_7_65, // sfix19_En18 
  input [18:0] Wgt_7_66, // sfix19_En18 
  input [18:0] Wgt_7_67, // sfix19_En18 
  input [18:0] Wgt_7_68, // sfix19_En18 
  input [18:0] Wgt_7_69, // sfix19_En18 
  input [18:0] Wgt_7_70, // sfix19_En18 
  input [18:0] Wgt_7_71, // sfix19_En18 
  input [18:0] Wgt_7_72, // sfix19_En18 
  input [18:0] Wgt_7_73, // sfix19_En18 
  input [18:0] Wgt_7_74, // sfix19_En18 
  input [18:0] Wgt_7_75, // sfix19_En18 
  input [18:0] Wgt_7_76, // sfix19_En18 
  input [18:0] Wgt_7_77, // sfix19_En18 
  input [18:0] Wgt_7_78, // sfix19_En18 
  input [18:0] Wgt_7_79, // sfix19_En18 
  input [18:0] Wgt_7_80, // sfix19_En18 
  input [18:0] Wgt_7_81, // sfix19_En18 
  input [18:0] Wgt_7_82, // sfix19_En18 
  input [18:0] Wgt_7_83, // sfix19_En18 
  input [18:0] Wgt_7_84, // sfix19_En18 
  input [18:0] Wgt_7_85, // sfix19_En18 
  input [18:0] Wgt_7_86, // sfix19_En18 
  input [18:0] Wgt_7_87, // sfix19_En18 
  input [18:0] Wgt_7_88, // sfix19_En18 
  input [18:0] Wgt_7_89, // sfix19_En18 
  input [18:0] Wgt_7_90, // sfix19_En18 
  input [18:0] Wgt_7_91, // sfix19_En18 
  input [18:0] Wgt_7_92, // sfix19_En18 
  input [18:0] Wgt_7_93, // sfix19_En18 
  input [18:0] Wgt_7_94, // sfix19_En18 
  input [18:0] Wgt_7_95, // sfix19_En18 
  input [18:0] Wgt_7_96, // sfix19_En18 
  input [18:0] Wgt_7_97, // sfix19_En18 
  input [18:0] Wgt_7_98, // sfix19_En18 
  input [18:0] Wgt_7_99, // sfix19_En18 
  input [18:0] Wgt_7_100, // sfix19_En18 
  input [18:0] Wgt_7_101, // sfix19_En18 
  input [18:0] Wgt_7_102, // sfix19_En18 
  input [18:0] Wgt_7_103, // sfix19_En18 
  input [18:0] Wgt_7_104, // sfix19_En18 
  input [18:0] Wgt_7_105, // sfix19_En18 
  input [18:0] Wgt_7_106, // sfix19_En18 
  input [18:0] Wgt_7_107, // sfix19_En18 
  input [18:0] Wgt_7_108, // sfix19_En18 
  input [18:0] Wgt_7_109, // sfix19_En18 
  input [18:0] Wgt_7_110, // sfix19_En18 
  input [18:0] Wgt_7_111, // sfix19_En18 
  input [18:0] Wgt_7_112, // sfix19_En18 
  input [18:0] Wgt_7_113, // sfix19_En18 
  input [18:0] Wgt_7_114, // sfix19_En18 
  input [18:0] Wgt_7_115, // sfix19_En18 
  input [18:0] Wgt_7_116, // sfix19_En18 
  input [18:0] Wgt_7_117, // sfix19_En18 
  input [18:0] Wgt_7_118, // sfix19_En18 
  input [18:0] Wgt_7_119, // sfix19_En18 
  input [18:0] Wgt_7_120, // sfix19_En18 
  input [18:0] Wgt_7_121, // sfix19_En18 
  input [18:0] Wgt_7_122, // sfix19_En18 
  input [18:0] Wgt_7_123, // sfix19_En18 
  input [18:0] Wgt_7_124, // sfix19_En18 
  input [18:0] Wgt_7_125, // sfix19_En18 
  input [18:0] Wgt_7_126, // sfix19_En18 
  input [18:0] Wgt_7_127, // sfix19_En18 
  input [18:0] Wgt_7_128, // sfix19_En18 
  input [18:0] Wgt_7_129, // sfix19_En18 
  input [18:0] Wgt_7_130, // sfix19_En18 
  input [18:0] Wgt_7_131, // sfix19_En18 
  input [18:0] Wgt_7_132, // sfix19_En18 
  input [18:0] Wgt_7_133, // sfix19_En18 
  input [18:0] Wgt_7_134, // sfix19_En18 
  input [18:0] Wgt_7_135, // sfix19_En18 
  input [18:0] Wgt_7_136, // sfix19_En18 
  input [18:0] Wgt_7_137, // sfix19_En18 
  input [18:0] Wgt_7_138, // sfix19_En18 
  input [18:0] Wgt_7_139, // sfix19_En18 
  input [18:0] Wgt_7_140, // sfix19_En18 
  input [18:0] Wgt_7_141, // sfix19_En18 
  input [18:0] Wgt_7_142, // sfix19_En18 
  input [18:0] Wgt_7_143, // sfix19_En18 
  input [18:0] Wgt_7_144, // sfix19_En18 
  input [18:0] Wgt_7_145, // sfix19_En18 
  input [18:0] Wgt_7_146, // sfix19_En18 
  input [18:0] Wgt_7_147, // sfix19_En18 
  input [18:0] Wgt_7_148, // sfix19_En18 
  input [18:0] Wgt_7_149, // sfix19_En18 
  input [18:0] Wgt_7_150, // sfix19_En18 
  input [18:0] Wgt_7_151, // sfix19_En18 
  input [18:0] Wgt_7_152, // sfix19_En18 
  input [18:0] Wgt_7_153, // sfix19_En18 
  input [18:0] Wgt_7_154, // sfix19_En18 
  input [18:0] Wgt_7_155, // sfix19_En18 
  input [18:0] Wgt_7_156, // sfix19_En18 
  input [18:0] Wgt_7_157, // sfix19_En18 
  input [18:0] Wgt_7_158, // sfix19_En18 
  input [18:0] Wgt_7_159, // sfix19_En18 
  input [18:0] Wgt_7_160, // sfix19_En18 
  input [18:0] Wgt_7_161, // sfix19_En18 
  input [18:0] Wgt_7_162, // sfix19_En18 
  input [18:0] Wgt_7_163, // sfix19_En18 
  input [18:0] Wgt_7_164, // sfix19_En18 
  input [18:0] Wgt_7_165, // sfix19_En18 
  input [18:0] Wgt_7_166, // sfix19_En18 
  input [18:0] Wgt_7_167, // sfix19_En18 
  input [18:0] Wgt_7_168, // sfix19_En18 
  input [18:0] Wgt_7_169, // sfix19_En18 
  input [18:0] Wgt_7_170, // sfix19_En18 
  input [18:0] Wgt_7_171, // sfix19_En18 
  input [18:0] Wgt_7_172, // sfix19_En18 
  input [18:0] Wgt_7_173, // sfix19_En18 
  input [18:0] Wgt_7_174, // sfix19_En18 
  input [18:0] Wgt_7_175, // sfix19_En18 
  input [18:0] Wgt_7_176, // sfix19_En18 
  input [18:0] Wgt_7_177, // sfix19_En18 
  input [18:0] Wgt_7_178, // sfix19_En18 
  input [18:0] Wgt_7_179, // sfix19_En18 
  input [18:0] Wgt_7_180, // sfix19_En18 
  input [18:0] Wgt_7_181, // sfix19_En18 
  input [18:0] Wgt_7_182, // sfix19_En18 
  input [18:0] Wgt_7_183, // sfix19_En18 
  input [18:0] Wgt_7_184, // sfix19_En18 
  input [18:0] Wgt_7_185, // sfix19_En18 
  input [18:0] Wgt_7_186, // sfix19_En18 
  input [18:0] Wgt_7_187, // sfix19_En18 
  input [18:0] Wgt_7_188, // sfix19_En18 
  input [18:0] Wgt_7_189, // sfix19_En18 
  input [18:0] Wgt_7_190, // sfix19_En18 
  input [18:0] Wgt_7_191, // sfix19_En18 
  input [18:0] Wgt_7_192, // sfix19_En18 
  input [18:0] Wgt_7_193, // sfix19_En18 
  input [18:0] Wgt_7_194, // sfix19_En18 
  input [18:0] Wgt_7_195, // sfix19_En18 
  input [18:0] Wgt_7_196, // sfix19_En18 
  input [18:0] Wgt_7_197, // sfix19_En18 
  input [18:0] Wgt_7_198, // sfix19_En18 
  input [18:0] Wgt_7_199, // sfix19_En18 
  input [18:0] Wgt_7_200, // sfix19_En18 
  input [18:0] Wgt_7_201, // sfix19_En18 
  input [18:0] Wgt_7_202, // sfix19_En18 
  input [18:0] Wgt_7_203, // sfix19_En18 
  input [18:0] Wgt_7_204, // sfix19_En18 
  input [18:0] Wgt_7_205, // sfix19_En18 
  input [18:0] Wgt_7_206, // sfix19_En18 
  input [18:0] Wgt_7_207, // sfix19_En18 
  input [18:0] Wgt_7_208, // sfix19_En18 
  input [18:0] Wgt_7_209, // sfix19_En18 
  input [18:0] Wgt_7_210, // sfix19_En18 
  input [18:0] Wgt_7_211, // sfix19_En18 
  input [18:0] Wgt_7_212, // sfix19_En18 
  input [18:0] Wgt_7_213, // sfix19_En18 
  input [18:0] Wgt_7_214, // sfix19_En18 
  input [18:0] Wgt_7_215, // sfix19_En18 
  input [18:0] Wgt_7_216, // sfix19_En18 
  input [18:0] Wgt_7_217, // sfix19_En18 
  input [18:0] Wgt_7_218, // sfix19_En18 
  input [18:0] Wgt_7_219, // sfix19_En18 
  input [18:0] Wgt_7_220, // sfix19_En18 
  input [18:0] Wgt_7_221, // sfix19_En18 
  input [18:0] Wgt_7_222, // sfix19_En18 
  input [18:0] Wgt_7_223, // sfix19_En18 
  input [18:0] Wgt_7_224, // sfix19_En18 
  input [18:0] Wgt_7_225, // sfix19_En18 
  input [18:0] Wgt_7_226, // sfix19_En18 
  input [18:0] Wgt_7_227, // sfix19_En18 
  input [18:0] Wgt_7_228, // sfix19_En18 
  input [18:0] Wgt_7_229, // sfix19_En18 
  input [18:0] Wgt_7_230, // sfix19_En18 
  input [18:0] Wgt_7_231, // sfix19_En18 
  input [18:0] Wgt_7_232, // sfix19_En18 
  input [18:0] Wgt_7_233, // sfix19_En18 
  input [18:0] Wgt_7_234, // sfix19_En18 
  input [18:0] Wgt_7_235, // sfix19_En18 
  input [18:0] Wgt_7_236, // sfix19_En18 
  input [18:0] Wgt_7_237, // sfix19_En18 
  input [18:0] Wgt_7_238, // sfix19_En18 
  input [18:0] Wgt_7_239, // sfix19_En18 
  input [18:0] Wgt_7_240, // sfix19_En18 
  input [18:0] Wgt_7_241, // sfix19_En18 
  input [18:0] Wgt_7_242, // sfix19_En18 
  input [18:0] Wgt_7_243, // sfix19_En18 
  input [18:0] Wgt_7_244, // sfix19_En18 
  input [18:0] Wgt_7_245, // sfix19_En18 
  input [18:0] Wgt_7_246, // sfix19_En18 
  input [18:0] Wgt_7_247, // sfix19_En18 
  input [18:0] Wgt_7_248, // sfix19_En18 
  input [18:0] Wgt_7_249, // sfix19_En18 
  input [18:0] Wgt_7_250, // sfix19_En18 
  input [18:0] Wgt_7_251, // sfix19_En18 
  input [18:0] Wgt_7_252, // sfix19_En18 
  input [18:0] Wgt_7_253, // sfix19_En18 
  input [18:0] Wgt_7_254, // sfix19_En18 
  input [18:0] Wgt_7_255, // sfix19_En18 
  input [18:0] Wgt_7_256, // sfix19_En18 
  input [18:0] Wgt_7_257, // sfix19_En18 
  input [18:0] Wgt_7_258, // sfix19_En18 
  input [18:0] Wgt_7_259, // sfix19_En18 
  input [18:0] Wgt_7_260, // sfix19_En18 
  input [18:0] Wgt_7_261, // sfix19_En18 
  input [18:0] Wgt_7_262, // sfix19_En18 
  input [18:0] Wgt_7_263, // sfix19_En18 
  input [18:0] Wgt_7_264, // sfix19_En18 
  input [18:0] Wgt_7_265, // sfix19_En18 
  input [18:0] Wgt_7_266, // sfix19_En18 
  input [18:0] Wgt_7_267, // sfix19_En18 
  input [18:0] Wgt_7_268, // sfix19_En18 
  input [18:0] Wgt_7_269, // sfix19_En18 
  input [18:0] Wgt_7_270, // sfix19_En18 
  input [18:0] Wgt_7_271, // sfix19_En18 
  input [18:0] Wgt_7_272, // sfix19_En18 
  input [18:0] Wgt_7_273, // sfix19_En18 
  input [18:0] Wgt_7_274, // sfix19_En18 
  input [18:0] Wgt_7_275, // sfix19_En18 
  input [18:0] Wgt_7_276, // sfix19_En18 
  input [18:0] Wgt_7_277, // sfix19_En18 
  input [18:0] Wgt_7_278, // sfix19_En18 
  input [18:0] Wgt_7_279, // sfix19_En18 
  input [18:0] Wgt_7_280, // sfix19_En18 
  input [18:0] Wgt_7_281, // sfix19_En18 
  input [18:0] Wgt_7_282, // sfix19_En18 
  input [18:0] Wgt_7_283, // sfix19_En18 
  input [18:0] Wgt_7_284, // sfix19_En18 
  input [18:0] Wgt_7_285, // sfix19_En18 
  input [18:0] Wgt_7_286, // sfix19_En18 
  input [18:0] Wgt_7_287, // sfix19_En18 
  input [18:0] Wgt_7_288, // sfix19_En18 
  input [18:0] Wgt_7_289, // sfix19_En18 
  input [18:0] Wgt_7_290, // sfix19_En18 
  input [18:0] Wgt_7_291, // sfix19_En18 
  input [18:0] Wgt_7_292, // sfix19_En18 
  input [18:0] Wgt_7_293, // sfix19_En18 
  input [18:0] Wgt_7_294, // sfix19_En18 
  input [18:0] Wgt_7_295, // sfix19_En18 
  input [18:0] Wgt_7_296, // sfix19_En18 
  input [18:0] Wgt_7_297, // sfix19_En18 
  input [18:0] Wgt_7_298, // sfix19_En18 
  input [18:0] Wgt_7_299, // sfix19_En18 
  input [18:0] Wgt_7_300, // sfix19_En18 
  input [18:0] Wgt_7_301, // sfix19_En18 
  input [18:0] Wgt_7_302, // sfix19_En18 
  input [18:0] Wgt_7_303, // sfix19_En18 
  input [18:0] Wgt_7_304, // sfix19_En18 
  input [18:0] Wgt_7_305, // sfix19_En18 
  input [18:0] Wgt_7_306, // sfix19_En18 
  input [18:0] Wgt_7_307, // sfix19_En18 
  input [18:0] Wgt_7_308, // sfix19_En18 
  input [18:0] Wgt_7_309, // sfix19_En18 
  input [18:0] Wgt_7_310, // sfix19_En18 
  input [18:0] Wgt_7_311, // sfix19_En18 
  input [18:0] Wgt_7_312, // sfix19_En18 
  input [18:0] Wgt_7_313, // sfix19_En18 
  input [18:0] Wgt_7_314, // sfix19_En18 
  input [18:0] Wgt_7_315, // sfix19_En18 
  input [18:0] Wgt_7_316, // sfix19_En18 
  input [18:0] Wgt_7_317, // sfix19_En18 
  input [18:0] Wgt_7_318, // sfix19_En18 
  input [18:0] Wgt_7_319, // sfix19_En18 
  input [18:0] Wgt_7_320, // sfix19_En18 
  input [18:0] Wgt_7_321, // sfix19_En18 
  input [18:0] Wgt_7_322, // sfix19_En18 
  input [18:0] Wgt_7_323, // sfix19_En18 
  input [18:0] Wgt_7_324, // sfix19_En18 
  input [18:0] Wgt_7_325, // sfix19_En18 
  input [18:0] Wgt_7_326, // sfix19_En18 
  input [18:0] Wgt_7_327, // sfix19_En18 
  input [18:0] Wgt_7_328, // sfix19_En18 
  input [18:0] Wgt_7_329, // sfix19_En18 
  input [18:0] Wgt_7_330, // sfix19_En18 
  input [18:0] Wgt_7_331, // sfix19_En18 
  input [18:0] Wgt_7_332, // sfix19_En18 
  input [18:0] Wgt_7_333, // sfix19_En18 
  input [18:0] Wgt_7_334, // sfix19_En18 
  input [18:0] Wgt_7_335, // sfix19_En18 
  input [18:0] Wgt_7_336, // sfix19_En18 
  input [18:0] Wgt_7_337, // sfix19_En18 
  input [18:0] Wgt_7_338, // sfix19_En18 
  input [18:0] Wgt_7_339, // sfix19_En18 
  input [18:0] Wgt_7_340, // sfix19_En18 
  input [18:0] Wgt_7_341, // sfix19_En18 
  input [18:0] Wgt_7_342, // sfix19_En18 
  input [18:0] Wgt_7_343, // sfix19_En18 
  input [18:0] Wgt_7_344, // sfix19_En18 
  input [18:0] Wgt_7_345, // sfix19_En18 
  input [18:0] Wgt_7_346, // sfix19_En18 
  input [18:0] Wgt_7_347, // sfix19_En18 
  input [18:0] Wgt_7_348, // sfix19_En18 
  input [18:0] Wgt_7_349, // sfix19_En18 
  input [18:0] Wgt_7_350, // sfix19_En18 
  input [18:0] Wgt_7_351, // sfix19_En18 
  input [18:0] Wgt_7_352, // sfix19_En18 
  input [18:0] Wgt_7_353, // sfix19_En18 
  input [18:0] Wgt_7_354, // sfix19_En18 
  input [18:0] Wgt_7_355, // sfix19_En18 
  input [18:0] Wgt_7_356, // sfix19_En18 
  input [18:0] Wgt_7_357, // sfix19_En18 
  input [18:0] Wgt_7_358, // sfix19_En18 
  input [18:0] Wgt_7_359, // sfix19_En18 
  input [18:0] Wgt_7_360, // sfix19_En18 
  input [18:0] Wgt_7_361, // sfix19_En18 
  input [18:0] Wgt_7_362, // sfix19_En18 
  input [18:0] Wgt_7_363, // sfix19_En18 
  input [18:0] Wgt_7_364, // sfix19_En18 
  input [18:0] Wgt_7_365, // sfix19_En18 
  input [18:0] Wgt_7_366, // sfix19_En18 
  input [18:0] Wgt_7_367, // sfix19_En18 
  input [18:0] Wgt_7_368, // sfix19_En18 
  input [18:0] Wgt_7_369, // sfix19_En18 
  input [18:0] Wgt_7_370, // sfix19_En18 
  input [18:0] Wgt_7_371, // sfix19_En18 
  input [18:0] Wgt_7_372, // sfix19_En18 
  input [18:0] Wgt_7_373, // sfix19_En18 
  input [18:0] Wgt_7_374, // sfix19_En18 
  input [18:0] Wgt_7_375, // sfix19_En18 
  input [18:0] Wgt_7_376, // sfix19_En18 
  input [18:0] Wgt_7_377, // sfix19_En18 
  input [18:0] Wgt_7_378, // sfix19_En18 
  input [18:0] Wgt_7_379, // sfix19_En18 
  input [18:0] Wgt_7_380, // sfix19_En18 
  input [18:0] Wgt_7_381, // sfix19_En18 
  input [18:0] Wgt_7_382, // sfix19_En18 
  input [18:0] Wgt_7_383, // sfix19_En18 
  input [18:0] Wgt_7_384, // sfix19_En18 
  input [18:0] Wgt_7_385, // sfix19_En18 
  input [18:0] Wgt_7_386, // sfix19_En18 
  input [18:0] Wgt_7_387, // sfix19_En18 
  input [18:0] Wgt_7_388, // sfix19_En18 
  input [18:0] Wgt_7_389, // sfix19_En18 
  input [18:0] Wgt_7_390, // sfix19_En18 
  input [18:0] Wgt_7_391, // sfix19_En18 
  input [18:0] Wgt_7_392, // sfix19_En18 
  input [18:0] Wgt_7_393, // sfix19_En18 
  input [18:0] Wgt_7_394, // sfix19_En18 
  input [18:0] Wgt_7_395, // sfix19_En18 
  input [18:0] Wgt_7_396, // sfix19_En18 
  input [18:0] Wgt_7_397, // sfix19_En18 
  input [18:0] Wgt_7_398, // sfix19_En18 
  input [18:0] Wgt_7_399, // sfix19_En18 
  input [18:0] Wgt_7_400, // sfix19_En18 
  input [18:0] Wgt_7_401, // sfix19_En18 
  input [18:0] Wgt_7_402, // sfix19_En18 
  input [18:0] Wgt_7_403, // sfix19_En18 
  input [18:0] Wgt_7_404, // sfix19_En18 
  input [18:0] Wgt_7_405, // sfix19_En18 
  input [18:0] Wgt_7_406, // sfix19_En18 
  input [18:0] Wgt_7_407, // sfix19_En18 
  input [18:0] Wgt_7_408, // sfix19_En18 
  input [18:0] Wgt_7_409, // sfix19_En18 
  input [18:0] Wgt_7_410, // sfix19_En18 
  input [18:0] Wgt_7_411, // sfix19_En18 
  input [18:0] Wgt_7_412, // sfix19_En18 
  input [18:0] Wgt_7_413, // sfix19_En18 
  input [18:0] Wgt_7_414, // sfix19_En18 
  input [18:0] Wgt_7_415, // sfix19_En18 
  input [18:0] Wgt_7_416, // sfix19_En18 
  input [18:0] Wgt_7_417, // sfix19_En18 
  input [18:0] Wgt_7_418, // sfix19_En18 
  input [18:0] Wgt_7_419, // sfix19_En18 
  input [18:0] Wgt_7_420, // sfix19_En18 
  input [18:0] Wgt_7_421, // sfix19_En18 
  input [18:0] Wgt_7_422, // sfix19_En18 
  input [18:0] Wgt_7_423, // sfix19_En18 
  input [18:0] Wgt_7_424, // sfix19_En18 
  input [18:0] Wgt_7_425, // sfix19_En18 
  input [18:0] Wgt_7_426, // sfix19_En18 
  input [18:0] Wgt_7_427, // sfix19_En18 
  input [18:0] Wgt_7_428, // sfix19_En18 
  input [18:0] Wgt_7_429, // sfix19_En18 
  input [18:0] Wgt_7_430, // sfix19_En18 
  input [18:0] Wgt_7_431, // sfix19_En18 
  input [18:0] Wgt_7_432, // sfix19_En18 
  input [18:0] Wgt_7_433, // sfix19_En18 
  input [18:0] Wgt_7_434, // sfix19_En18 
  input [18:0] Wgt_7_435, // sfix19_En18 
  input [18:0] Wgt_7_436, // sfix19_En18 
  input [18:0] Wgt_7_437, // sfix19_En18 
  input [18:0] Wgt_7_438, // sfix19_En18 
  input [18:0] Wgt_7_439, // sfix19_En18 
  input [18:0] Wgt_7_440, // sfix19_En18 
  input [18:0] Wgt_7_441, // sfix19_En18 
  input [18:0] Wgt_7_442, // sfix19_En18 
  input [18:0] Wgt_7_443, // sfix19_En18 
  input [18:0] Wgt_7_444, // sfix19_En18 
  input [18:0] Wgt_7_445, // sfix19_En18 
  input [18:0] Wgt_7_446, // sfix19_En18 
  input [18:0] Wgt_7_447, // sfix19_En18 
  input [18:0] Wgt_7_448, // sfix19_En18 
  input [18:0] Wgt_7_449, // sfix19_En18 
  input [18:0] Wgt_7_450, // sfix19_En18 
  input [18:0] Wgt_7_451, // sfix19_En18 
  input [18:0] Wgt_7_452, // sfix19_En18 
  input [18:0] Wgt_7_453, // sfix19_En18 
  input [18:0] Wgt_7_454, // sfix19_En18 
  input [18:0] Wgt_7_455, // sfix19_En18 
  input [18:0] Wgt_7_456, // sfix19_En18 
  input [18:0] Wgt_7_457, // sfix19_En18 
  input [18:0] Wgt_7_458, // sfix19_En18 
  input [18:0] Wgt_7_459, // sfix19_En18 
  input [18:0] Wgt_7_460, // sfix19_En18 
  input [18:0] Wgt_7_461, // sfix19_En18 
  input [18:0] Wgt_7_462, // sfix19_En18 
  input [18:0] Wgt_7_463, // sfix19_En18 
  input [18:0] Wgt_7_464, // sfix19_En18 
  input [18:0] Wgt_7_465, // sfix19_En18 
  input [18:0] Wgt_7_466, // sfix19_En18 
  input [18:0] Wgt_7_467, // sfix19_En18 
  input [18:0] Wgt_7_468, // sfix19_En18 
  input [18:0] Wgt_7_469, // sfix19_En18 
  input [18:0] Wgt_7_470, // sfix19_En18 
  input [18:0] Wgt_7_471, // sfix19_En18 
  input [18:0] Wgt_7_472, // sfix19_En18 
  input [18:0] Wgt_7_473, // sfix19_En18 
  input [18:0] Wgt_7_474, // sfix19_En18 
  input [18:0] Wgt_7_475, // sfix19_En18 
  input [18:0] Wgt_7_476, // sfix19_En18 
  input [18:0] Wgt_7_477, // sfix19_En18 
  input [18:0] Wgt_7_478, // sfix19_En18 
  input [18:0] Wgt_7_479, // sfix19_En18 
  input [18:0] Wgt_7_480, // sfix19_En18 
  input [18:0] Wgt_7_481, // sfix19_En18 
  input [18:0] Wgt_7_482, // sfix19_En18 
  input [18:0] Wgt_7_483, // sfix19_En18 
  input [18:0] Wgt_7_484, // sfix19_En18 
  input [18:0] Wgt_7_485, // sfix19_En18 
  input [18:0] Wgt_7_486, // sfix19_En18 
  input [18:0] Wgt_7_487, // sfix19_En18 
  input [18:0] Wgt_7_488, // sfix19_En18 
  input [18:0] Wgt_7_489, // sfix19_En18 
  input [18:0] Wgt_7_490, // sfix19_En18 
  input [18:0] Wgt_7_491, // sfix19_En18 
  input [18:0] Wgt_7_492, // sfix19_En18 
  input [18:0] Wgt_7_493, // sfix19_En18 
  input [18:0] Wgt_7_494, // sfix19_En18 
  input [18:0] Wgt_7_495, // sfix19_En18 
  input [18:0] Wgt_7_496, // sfix19_En18 
  input [18:0] Wgt_7_497, // sfix19_En18 
  input [18:0] Wgt_7_498, // sfix19_En18 
  input [18:0] Wgt_7_499, // sfix19_En18 
  input [18:0] Wgt_7_500, // sfix19_En18 
  input [18:0] Wgt_7_501, // sfix19_En18 
  input [18:0] Wgt_7_502, // sfix19_En18 
  input [18:0] Wgt_7_503, // sfix19_En18 
  input [18:0] Wgt_7_504, // sfix19_En18 
  input [18:0] Wgt_7_505, // sfix19_En18 
  input [18:0] Wgt_7_506, // sfix19_En18 
  input [18:0] Wgt_7_507, // sfix19_En18 
  input [18:0] Wgt_7_508, // sfix19_En18 
  input [18:0] Wgt_7_509, // sfix19_En18 
  input [18:0] Wgt_7_510, // sfix19_En18 
  input [18:0] Wgt_7_511, // sfix19_En18 
  input [18:0] Wgt_7_512, // sfix19_En18 
  input [18:0] Wgt_7_513, // sfix19_En18 
  input [18:0] Wgt_7_514, // sfix19_En18 
  input [18:0] Wgt_7_515, // sfix19_En18 
  input [18:0] Wgt_7_516, // sfix19_En18 
  input [18:0] Wgt_7_517, // sfix19_En18 
  input [18:0] Wgt_7_518, // sfix19_En18 
  input [18:0] Wgt_7_519, // sfix19_En18 
  input [18:0] Wgt_7_520, // sfix19_En18 
  input [18:0] Wgt_7_521, // sfix19_En18 
  input [18:0] Wgt_7_522, // sfix19_En18 
  input [18:0] Wgt_7_523, // sfix19_En18 
  input [18:0] Wgt_7_524, // sfix19_En18 
  input [18:0] Wgt_7_525, // sfix19_En18 
  input [18:0] Wgt_7_526, // sfix19_En18 
  input [18:0] Wgt_7_527, // sfix19_En18 
  input [18:0] Wgt_7_528, // sfix19_En18 
  input [18:0] Wgt_7_529, // sfix19_En18 
  input [18:0] Wgt_7_530, // sfix19_En18 
  input [18:0] Wgt_7_531, // sfix19_En18 
  input [18:0] Wgt_7_532, // sfix19_En18 
  input [18:0] Wgt_7_533, // sfix19_En18 
  input [18:0] Wgt_7_534, // sfix19_En18 
  input [18:0] Wgt_7_535, // sfix19_En18 
  input [18:0] Wgt_7_536, // sfix19_En18 
  input [18:0] Wgt_7_537, // sfix19_En18 
  input [18:0] Wgt_7_538, // sfix19_En18 
  input [18:0] Wgt_7_539, // sfix19_En18 
  input [18:0] Wgt_7_540, // sfix19_En18 
  input [18:0] Wgt_7_541, // sfix19_En18 
  input [18:0] Wgt_7_542, // sfix19_En18 
  input [18:0] Wgt_7_543, // sfix19_En18 
  input [18:0] Wgt_7_544, // sfix19_En18 
  input [18:0] Wgt_7_545, // sfix19_En18 
  input [18:0] Wgt_7_546, // sfix19_En18 
  input [18:0] Wgt_7_547, // sfix19_En18 
  input [18:0] Wgt_7_548, // sfix19_En18 
  input [18:0] Wgt_7_549, // sfix19_En18 
  input [18:0] Wgt_7_550, // sfix19_En18 
  input [18:0] Wgt_7_551, // sfix19_En18 
  input [18:0] Wgt_7_552, // sfix19_En18 
  input [18:0] Wgt_7_553, // sfix19_En18 
  input [18:0] Wgt_7_554, // sfix19_En18 
  input [18:0] Wgt_7_555, // sfix19_En18 
  input [18:0] Wgt_7_556, // sfix19_En18 
  input [18:0] Wgt_7_557, // sfix19_En18 
  input [18:0] Wgt_7_558, // sfix19_En18 
  input [18:0] Wgt_7_559, // sfix19_En18 
  input [18:0] Wgt_7_560, // sfix19_En18 
  input [18:0] Wgt_7_561, // sfix19_En18 
  input [18:0] Wgt_7_562, // sfix19_En18 
  input [18:0] Wgt_7_563, // sfix19_En18 
  input [18:0] Wgt_7_564, // sfix19_En18 
  input [18:0] Wgt_7_565, // sfix19_En18 
  input [18:0] Wgt_7_566, // sfix19_En18 
  input [18:0] Wgt_7_567, // sfix19_En18 
  input [18:0] Wgt_7_568, // sfix19_En18 
  input [18:0] Wgt_7_569, // sfix19_En18 
  input [18:0] Wgt_7_570, // sfix19_En18 
  input [18:0] Wgt_7_571, // sfix19_En18 
  input [18:0] Wgt_7_572, // sfix19_En18 
  input [18:0] Wgt_7_573, // sfix19_En18 
  input [18:0] Wgt_7_574, // sfix19_En18 
  input [18:0] Wgt_7_575, // sfix19_En18 
  input [18:0] Wgt_7_576, // sfix19_En18 
  input [18:0] Wgt_7_577, // sfix19_En18 
  input [18:0] Wgt_7_578, // sfix19_En18 
  input [18:0] Wgt_7_579, // sfix19_En18 
  input [18:0] Wgt_7_580, // sfix19_En18 
  input [18:0] Wgt_7_581, // sfix19_En18 
  input [18:0] Wgt_7_582, // sfix19_En18 
  input [18:0] Wgt_7_583, // sfix19_En18 
  input [18:0] Wgt_7_584, // sfix19_En18 
  input [18:0] Wgt_7_585, // sfix19_En18 
  input [18:0] Wgt_7_586, // sfix19_En18 
  input [18:0] Wgt_7_587, // sfix19_En18 
  input [18:0] Wgt_7_588, // sfix19_En18 
  input [18:0] Wgt_7_589, // sfix19_En18 
  input [18:0] Wgt_7_590, // sfix19_En18 
  input [18:0] Wgt_7_591, // sfix19_En18 
  input [18:0] Wgt_7_592, // sfix19_En18 
  input [18:0] Wgt_7_593, // sfix19_En18 
  input [18:0] Wgt_7_594, // sfix19_En18 
  input [18:0] Wgt_7_595, // sfix19_En18 
  input [18:0] Wgt_7_596, // sfix19_En18 
  input [18:0] Wgt_7_597, // sfix19_En18 
  input [18:0] Wgt_7_598, // sfix19_En18 
  input [18:0] Wgt_7_599, // sfix19_En18 
  input [18:0] Wgt_7_600, // sfix19_En18 
  input [18:0] Wgt_7_601, // sfix19_En18 
  input [18:0] Wgt_7_602, // sfix19_En18 
  input [18:0] Wgt_7_603, // sfix19_En18 
  input [18:0] Wgt_7_604, // sfix19_En18 
  input [18:0] Wgt_7_605, // sfix19_En18 
  input [18:0] Wgt_7_606, // sfix19_En18 
  input [18:0] Wgt_7_607, // sfix19_En18 
  input [18:0] Wgt_7_608, // sfix19_En18 
  input [18:0] Wgt_7_609, // sfix19_En18 
  input [18:0] Wgt_7_610, // sfix19_En18 
  input [18:0] Wgt_7_611, // sfix19_En18 
  input [18:0] Wgt_7_612, // sfix19_En18 
  input [18:0] Wgt_7_613, // sfix19_En18 
  input [18:0] Wgt_7_614, // sfix19_En18 
  input [18:0] Wgt_7_615, // sfix19_En18 
  input [18:0] Wgt_7_616, // sfix19_En18 
  input [18:0] Wgt_7_617, // sfix19_En18 
  input [18:0] Wgt_7_618, // sfix19_En18 
  input [18:0] Wgt_7_619, // sfix19_En18 
  input [18:0] Wgt_7_620, // sfix19_En18 
  input [18:0] Wgt_7_621, // sfix19_En18 
  input [18:0] Wgt_7_622, // sfix19_En18 
  input [18:0] Wgt_7_623, // sfix19_En18 
  input [18:0] Wgt_7_624, // sfix19_En18 
  input [18:0] Wgt_7_625, // sfix19_En18 
  input [18:0] Wgt_7_626, // sfix19_En18 
  input [18:0] Wgt_7_627, // sfix19_En18 
  input [18:0] Wgt_7_628, // sfix19_En18 
  input [18:0] Wgt_7_629, // sfix19_En18 
  input [18:0] Wgt_7_630, // sfix19_En18 
  input [18:0] Wgt_7_631, // sfix19_En18 
  input [18:0] Wgt_7_632, // sfix19_En18 
  input [18:0] Wgt_7_633, // sfix19_En18 
  input [18:0] Wgt_7_634, // sfix19_En18 
  input [18:0] Wgt_7_635, // sfix19_En18 
  input [18:0] Wgt_7_636, // sfix19_En18 
  input [18:0] Wgt_7_637, // sfix19_En18 
  input [18:0] Wgt_7_638, // sfix19_En18 
  input [18:0] Wgt_7_639, // sfix19_En18 
  input [18:0] Wgt_7_640, // sfix19_En18 
  input [18:0] Wgt_7_641, // sfix19_En18 
  input [18:0] Wgt_7_642, // sfix19_En18 
  input [18:0] Wgt_7_643, // sfix19_En18 
  input [18:0] Wgt_7_644, // sfix19_En18 
  input [18:0] Wgt_7_645, // sfix19_En18 
  input [18:0] Wgt_7_646, // sfix19_En18 
  input [18:0] Wgt_7_647, // sfix19_En18 
  input [18:0] Wgt_7_648, // sfix19_En18 
  input [18:0] Wgt_7_649, // sfix19_En18 
  input [18:0] Wgt_7_650, // sfix19_En18 
  input [18:0] Wgt_7_651, // sfix19_En18 
  input [18:0] Wgt_7_652, // sfix19_En18 
  input [18:0] Wgt_7_653, // sfix19_En18 
  input [18:0] Wgt_7_654, // sfix19_En18 
  input [18:0] Wgt_7_655, // sfix19_En18 
  input [18:0] Wgt_7_656, // sfix19_En18 
  input [18:0] Wgt_7_657, // sfix19_En18 
  input [18:0] Wgt_7_658, // sfix19_En18 
  input [18:0] Wgt_7_659, // sfix19_En18 
  input [18:0] Wgt_7_660, // sfix19_En18 
  input [18:0] Wgt_7_661, // sfix19_En18 
  input [18:0] Wgt_7_662, // sfix19_En18 
  input [18:0] Wgt_7_663, // sfix19_En18 
  input [18:0] Wgt_7_664, // sfix19_En18 
  input [18:0] Wgt_7_665, // sfix19_En18 
  input [18:0] Wgt_7_666, // sfix19_En18 
  input [18:0] Wgt_7_667, // sfix19_En18 
  input [18:0] Wgt_7_668, // sfix19_En18 
  input [18:0] Wgt_7_669, // sfix19_En18 
  input [18:0] Wgt_7_670, // sfix19_En18 
  input [18:0] Wgt_7_671, // sfix19_En18 
  input [18:0] Wgt_7_672, // sfix19_En18 
  input [18:0] Wgt_7_673, // sfix19_En18 
  input [18:0] Wgt_7_674, // sfix19_En18 
  input [18:0] Wgt_7_675, // sfix19_En18 
  input [18:0] Wgt_7_676, // sfix19_En18 
  input [18:0] Wgt_7_677, // sfix19_En18 
  input [18:0] Wgt_7_678, // sfix19_En18 
  input [18:0] Wgt_7_679, // sfix19_En18 
  input [18:0] Wgt_7_680, // sfix19_En18 
  input [18:0] Wgt_7_681, // sfix19_En18 
  input [18:0] Wgt_7_682, // sfix19_En18 
  input [18:0] Wgt_7_683, // sfix19_En18 
  input [18:0] Wgt_7_684, // sfix19_En18 
  input [18:0] Wgt_7_685, // sfix19_En18 
  input [18:0] Wgt_7_686, // sfix19_En18 
  input [18:0] Wgt_7_687, // sfix19_En18 
  input [18:0] Wgt_7_688, // sfix19_En18 
  input [18:0] Wgt_7_689, // sfix19_En18 
  input [18:0] Wgt_7_690, // sfix19_En18 
  input [18:0] Wgt_7_691, // sfix19_En18 
  input [18:0] Wgt_7_692, // sfix19_En18 
  input [18:0] Wgt_7_693, // sfix19_En18 
  input [18:0] Wgt_7_694, // sfix19_En18 
  input [18:0] Wgt_7_695, // sfix19_En18 
  input [18:0] Wgt_7_696, // sfix19_En18 
  input [18:0] Wgt_7_697, // sfix19_En18 
  input [18:0] Wgt_7_698, // sfix19_En18 
  input [18:0] Wgt_7_699, // sfix19_En18 
  input [18:0] Wgt_7_700, // sfix19_En18 
  input [18:0] Wgt_7_701, // sfix19_En18 
  input [18:0] Wgt_7_702, // sfix19_En18 
  input [18:0] Wgt_7_703, // sfix19_En18 
  input [18:0] Wgt_7_704, // sfix19_En18 
  input [18:0] Wgt_7_705, // sfix19_En18 
  input [18:0] Wgt_7_706, // sfix19_En18 
  input [18:0] Wgt_7_707, // sfix19_En18 
  input [18:0] Wgt_7_708, // sfix19_En18 
  input [18:0] Wgt_7_709, // sfix19_En18 
  input [18:0] Wgt_7_710, // sfix19_En18 
  input [18:0] Wgt_7_711, // sfix19_En18 
  input [18:0] Wgt_7_712, // sfix19_En18 
  input [18:0] Wgt_7_713, // sfix19_En18 
  input [18:0] Wgt_7_714, // sfix19_En18 
  input [18:0] Wgt_7_715, // sfix19_En18 
  input [18:0] Wgt_7_716, // sfix19_En18 
  input [18:0] Wgt_7_717, // sfix19_En18 
  input [18:0] Wgt_7_718, // sfix19_En18 
  input [18:0] Wgt_7_719, // sfix19_En18 
  input [18:0] Wgt_7_720, // sfix19_En18 
  input [18:0] Wgt_7_721, // sfix19_En18 
  input [18:0] Wgt_7_722, // sfix19_En18 
  input [18:0] Wgt_7_723, // sfix19_En18 
  input [18:0] Wgt_7_724, // sfix19_En18 
  input [18:0] Wgt_7_725, // sfix19_En18 
  input [18:0] Wgt_7_726, // sfix19_En18 
  input [18:0] Wgt_7_727, // sfix19_En18 
  input [18:0] Wgt_7_728, // sfix19_En18 
  input [18:0] Wgt_7_729, // sfix19_En18 
  input [18:0] Wgt_7_730, // sfix19_En18 
  input [18:0] Wgt_7_731, // sfix19_En18 
  input [18:0] Wgt_7_732, // sfix19_En18 
  input [18:0] Wgt_7_733, // sfix19_En18 
  input [18:0] Wgt_7_734, // sfix19_En18 
  input [18:0] Wgt_7_735, // sfix19_En18 
  input [18:0] Wgt_7_736, // sfix19_En18 
  input [18:0] Wgt_7_737, // sfix19_En18 
  input [18:0] Wgt_7_738, // sfix19_En18 
  input [18:0] Wgt_7_739, // sfix19_En18 
  input [18:0] Wgt_7_740, // sfix19_En18 
  input [18:0] Wgt_7_741, // sfix19_En18 
  input [18:0] Wgt_7_742, // sfix19_En18 
  input [18:0] Wgt_7_743, // sfix19_En18 
  input [18:0] Wgt_7_744, // sfix19_En18 
  input [18:0] Wgt_7_745, // sfix19_En18 
  input [18:0] Wgt_7_746, // sfix19_En18 
  input [18:0] Wgt_7_747, // sfix19_En18 
  input [18:0] Wgt_7_748, // sfix19_En18 
  input [18:0] Wgt_7_749, // sfix19_En18 
  input [18:0] Wgt_7_750, // sfix19_En18 
  input [18:0] Wgt_7_751, // sfix19_En18 
  input [18:0] Wgt_7_752, // sfix19_En18 
  input [18:0] Wgt_7_753, // sfix19_En18 
  input [18:0] Wgt_7_754, // sfix19_En18 
  input [18:0] Wgt_7_755, // sfix19_En18 
  input [18:0] Wgt_7_756, // sfix19_En18 
  input [18:0] Wgt_7_757, // sfix19_En18 
  input [18:0] Wgt_7_758, // sfix19_En18 
  input [18:0] Wgt_7_759, // sfix19_En18 
  input [18:0] Wgt_7_760, // sfix19_En18 
  input [18:0] Wgt_7_761, // sfix19_En18 
  input [18:0] Wgt_7_762, // sfix19_En18 
  input [18:0] Wgt_7_763, // sfix19_En18 
  input [18:0] Wgt_7_764, // sfix19_En18 
  input [18:0] Wgt_7_765, // sfix19_En18 
  input [18:0] Wgt_7_766, // sfix19_En18 
  input [18:0] Wgt_7_767, // sfix19_En18 
  input [18:0] Wgt_7_768, // sfix19_En18 
  input [18:0] Wgt_7_769, // sfix19_En18 
  input [18:0] Wgt_7_770, // sfix19_En18 
  input [18:0] Wgt_7_771, // sfix19_En18 
  input [18:0] Wgt_7_772, // sfix19_En18 
  input [18:0] Wgt_7_773, // sfix19_En18 
  input [18:0] Wgt_7_774, // sfix19_En18 
  input [18:0] Wgt_7_775, // sfix19_En18 
  input [18:0] Wgt_7_776, // sfix19_En18 
  input [18:0] Wgt_7_777, // sfix19_En18 
  input [18:0] Wgt_7_778, // sfix19_En18 
  input [18:0] Wgt_7_779, // sfix19_En18 
  input [18:0] Wgt_7_780, // sfix19_En18 
  input [18:0] Wgt_7_781, // sfix19_En18 
  input [18:0] Wgt_7_782, // sfix19_En18 
  input [18:0] Wgt_7_783, // sfix19_En18 
  input [18:0] Wgt_7_784, // sfix19_En18 
  input [18:0] Wgt_8_0, // sfix19_En18 
  input [18:0] Wgt_8_1, // sfix19_En18 
  input [18:0] Wgt_8_2, // sfix19_En18 
  input [18:0] Wgt_8_3, // sfix19_En18 
  input [18:0] Wgt_8_4, // sfix19_En18 
  input [18:0] Wgt_8_5, // sfix19_En18 
  input [18:0] Wgt_8_6, // sfix19_En18 
  input [18:0] Wgt_8_7, // sfix19_En18 
  input [18:0] Wgt_8_8, // sfix19_En18 
  input [18:0] Wgt_8_9, // sfix19_En18 
  input [18:0] Wgt_8_10, // sfix19_En18 
  input [18:0] Wgt_8_11, // sfix19_En18 
  input [18:0] Wgt_8_12, // sfix19_En18 
  input [18:0] Wgt_8_13, // sfix19_En18 
  input [18:0] Wgt_8_14, // sfix19_En18 
  input [18:0] Wgt_8_15, // sfix19_En18 
  input [18:0] Wgt_8_16, // sfix19_En18 
  input [18:0] Wgt_8_17, // sfix19_En18 
  input [18:0] Wgt_8_18, // sfix19_En18 
  input [18:0] Wgt_8_19, // sfix19_En18 
  input [18:0] Wgt_8_20, // sfix19_En18 
  input [18:0] Wgt_8_21, // sfix19_En18 
  input [18:0] Wgt_8_22, // sfix19_En18 
  input [18:0] Wgt_8_23, // sfix19_En18 
  input [18:0] Wgt_8_24, // sfix19_En18 
  input [18:0] Wgt_8_25, // sfix19_En18 
  input [18:0] Wgt_8_26, // sfix19_En18 
  input [18:0] Wgt_8_27, // sfix19_En18 
  input [18:0] Wgt_8_28, // sfix19_En18 
  input [18:0] Wgt_8_29, // sfix19_En18 
  input [18:0] Wgt_8_30, // sfix19_En18 
  input [18:0] Wgt_8_31, // sfix19_En18 
  input [18:0] Wgt_8_32, // sfix19_En18 
  input [18:0] Wgt_8_33, // sfix19_En18 
  input [18:0] Wgt_8_34, // sfix19_En18 
  input [18:0] Wgt_8_35, // sfix19_En18 
  input [18:0] Wgt_8_36, // sfix19_En18 
  input [18:0] Wgt_8_37, // sfix19_En18 
  input [18:0] Wgt_8_38, // sfix19_En18 
  input [18:0] Wgt_8_39, // sfix19_En18 
  input [18:0] Wgt_8_40, // sfix19_En18 
  input [18:0] Wgt_8_41, // sfix19_En18 
  input [18:0] Wgt_8_42, // sfix19_En18 
  input [18:0] Wgt_8_43, // sfix19_En18 
  input [18:0] Wgt_8_44, // sfix19_En18 
  input [18:0] Wgt_8_45, // sfix19_En18 
  input [18:0] Wgt_8_46, // sfix19_En18 
  input [18:0] Wgt_8_47, // sfix19_En18 
  input [18:0] Wgt_8_48, // sfix19_En18 
  input [18:0] Wgt_8_49, // sfix19_En18 
  input [18:0] Wgt_8_50, // sfix19_En18 
  input [18:0] Wgt_8_51, // sfix19_En18 
  input [18:0] Wgt_8_52, // sfix19_En18 
  input [18:0] Wgt_8_53, // sfix19_En18 
  input [18:0] Wgt_8_54, // sfix19_En18 
  input [18:0] Wgt_8_55, // sfix19_En18 
  input [18:0] Wgt_8_56, // sfix19_En18 
  input [18:0] Wgt_8_57, // sfix19_En18 
  input [18:0] Wgt_8_58, // sfix19_En18 
  input [18:0] Wgt_8_59, // sfix19_En18 
  input [18:0] Wgt_8_60, // sfix19_En18 
  input [18:0] Wgt_8_61, // sfix19_En18 
  input [18:0] Wgt_8_62, // sfix19_En18 
  input [18:0] Wgt_8_63, // sfix19_En18 
  input [18:0] Wgt_8_64, // sfix19_En18 
  input [18:0] Wgt_8_65, // sfix19_En18 
  input [18:0] Wgt_8_66, // sfix19_En18 
  input [18:0] Wgt_8_67, // sfix19_En18 
  input [18:0] Wgt_8_68, // sfix19_En18 
  input [18:0] Wgt_8_69, // sfix19_En18 
  input [18:0] Wgt_8_70, // sfix19_En18 
  input [18:0] Wgt_8_71, // sfix19_En18 
  input [18:0] Wgt_8_72, // sfix19_En18 
  input [18:0] Wgt_8_73, // sfix19_En18 
  input [18:0] Wgt_8_74, // sfix19_En18 
  input [18:0] Wgt_8_75, // sfix19_En18 
  input [18:0] Wgt_8_76, // sfix19_En18 
  input [18:0] Wgt_8_77, // sfix19_En18 
  input [18:0] Wgt_8_78, // sfix19_En18 
  input [18:0] Wgt_8_79, // sfix19_En18 
  input [18:0] Wgt_8_80, // sfix19_En18 
  input [18:0] Wgt_8_81, // sfix19_En18 
  input [18:0] Wgt_8_82, // sfix19_En18 
  input [18:0] Wgt_8_83, // sfix19_En18 
  input [18:0] Wgt_8_84, // sfix19_En18 
  input [18:0] Wgt_8_85, // sfix19_En18 
  input [18:0] Wgt_8_86, // sfix19_En18 
  input [18:0] Wgt_8_87, // sfix19_En18 
  input [18:0] Wgt_8_88, // sfix19_En18 
  input [18:0] Wgt_8_89, // sfix19_En18 
  input [18:0] Wgt_8_90, // sfix19_En18 
  input [18:0] Wgt_8_91, // sfix19_En18 
  input [18:0] Wgt_8_92, // sfix19_En18 
  input [18:0] Wgt_8_93, // sfix19_En18 
  input [18:0] Wgt_8_94, // sfix19_En18 
  input [18:0] Wgt_8_95, // sfix19_En18 
  input [18:0] Wgt_8_96, // sfix19_En18 
  input [18:0] Wgt_8_97, // sfix19_En18 
  input [18:0] Wgt_8_98, // sfix19_En18 
  input [18:0] Wgt_8_99, // sfix19_En18 
  input [18:0] Wgt_8_100, // sfix19_En18 
  input [18:0] Wgt_8_101, // sfix19_En18 
  input [18:0] Wgt_8_102, // sfix19_En18 
  input [18:0] Wgt_8_103, // sfix19_En18 
  input [18:0] Wgt_8_104, // sfix19_En18 
  input [18:0] Wgt_8_105, // sfix19_En18 
  input [18:0] Wgt_8_106, // sfix19_En18 
  input [18:0] Wgt_8_107, // sfix19_En18 
  input [18:0] Wgt_8_108, // sfix19_En18 
  input [18:0] Wgt_8_109, // sfix19_En18 
  input [18:0] Wgt_8_110, // sfix19_En18 
  input [18:0] Wgt_8_111, // sfix19_En18 
  input [18:0] Wgt_8_112, // sfix19_En18 
  input [18:0] Wgt_8_113, // sfix19_En18 
  input [18:0] Wgt_8_114, // sfix19_En18 
  input [18:0] Wgt_8_115, // sfix19_En18 
  input [18:0] Wgt_8_116, // sfix19_En18 
  input [18:0] Wgt_8_117, // sfix19_En18 
  input [18:0] Wgt_8_118, // sfix19_En18 
  input [18:0] Wgt_8_119, // sfix19_En18 
  input [18:0] Wgt_8_120, // sfix19_En18 
  input [18:0] Wgt_8_121, // sfix19_En18 
  input [18:0] Wgt_8_122, // sfix19_En18 
  input [18:0] Wgt_8_123, // sfix19_En18 
  input [18:0] Wgt_8_124, // sfix19_En18 
  input [18:0] Wgt_8_125, // sfix19_En18 
  input [18:0] Wgt_8_126, // sfix19_En18 
  input [18:0] Wgt_8_127, // sfix19_En18 
  input [18:0] Wgt_8_128, // sfix19_En18 
  input [18:0] Wgt_8_129, // sfix19_En18 
  input [18:0] Wgt_8_130, // sfix19_En18 
  input [18:0] Wgt_8_131, // sfix19_En18 
  input [18:0] Wgt_8_132, // sfix19_En18 
  input [18:0] Wgt_8_133, // sfix19_En18 
  input [18:0] Wgt_8_134, // sfix19_En18 
  input [18:0] Wgt_8_135, // sfix19_En18 
  input [18:0] Wgt_8_136, // sfix19_En18 
  input [18:0] Wgt_8_137, // sfix19_En18 
  input [18:0] Wgt_8_138, // sfix19_En18 
  input [18:0] Wgt_8_139, // sfix19_En18 
  input [18:0] Wgt_8_140, // sfix19_En18 
  input [18:0] Wgt_8_141, // sfix19_En18 
  input [18:0] Wgt_8_142, // sfix19_En18 
  input [18:0] Wgt_8_143, // sfix19_En18 
  input [18:0] Wgt_8_144, // sfix19_En18 
  input [18:0] Wgt_8_145, // sfix19_En18 
  input [18:0] Wgt_8_146, // sfix19_En18 
  input [18:0] Wgt_8_147, // sfix19_En18 
  input [18:0] Wgt_8_148, // sfix19_En18 
  input [18:0] Wgt_8_149, // sfix19_En18 
  input [18:0] Wgt_8_150, // sfix19_En18 
  input [18:0] Wgt_8_151, // sfix19_En18 
  input [18:0] Wgt_8_152, // sfix19_En18 
  input [18:0] Wgt_8_153, // sfix19_En18 
  input [18:0] Wgt_8_154, // sfix19_En18 
  input [18:0] Wgt_8_155, // sfix19_En18 
  input [18:0] Wgt_8_156, // sfix19_En18 
  input [18:0] Wgt_8_157, // sfix19_En18 
  input [18:0] Wgt_8_158, // sfix19_En18 
  input [18:0] Wgt_8_159, // sfix19_En18 
  input [18:0] Wgt_8_160, // sfix19_En18 
  input [18:0] Wgt_8_161, // sfix19_En18 
  input [18:0] Wgt_8_162, // sfix19_En18 
  input [18:0] Wgt_8_163, // sfix19_En18 
  input [18:0] Wgt_8_164, // sfix19_En18 
  input [18:0] Wgt_8_165, // sfix19_En18 
  input [18:0] Wgt_8_166, // sfix19_En18 
  input [18:0] Wgt_8_167, // sfix19_En18 
  input [18:0] Wgt_8_168, // sfix19_En18 
  input [18:0] Wgt_8_169, // sfix19_En18 
  input [18:0] Wgt_8_170, // sfix19_En18 
  input [18:0] Wgt_8_171, // sfix19_En18 
  input [18:0] Wgt_8_172, // sfix19_En18 
  input [18:0] Wgt_8_173, // sfix19_En18 
  input [18:0] Wgt_8_174, // sfix19_En18 
  input [18:0] Wgt_8_175, // sfix19_En18 
  input [18:0] Wgt_8_176, // sfix19_En18 
  input [18:0] Wgt_8_177, // sfix19_En18 
  input [18:0] Wgt_8_178, // sfix19_En18 
  input [18:0] Wgt_8_179, // sfix19_En18 
  input [18:0] Wgt_8_180, // sfix19_En18 
  input [18:0] Wgt_8_181, // sfix19_En18 
  input [18:0] Wgt_8_182, // sfix19_En18 
  input [18:0] Wgt_8_183, // sfix19_En18 
  input [18:0] Wgt_8_184, // sfix19_En18 
  input [18:0] Wgt_8_185, // sfix19_En18 
  input [18:0] Wgt_8_186, // sfix19_En18 
  input [18:0] Wgt_8_187, // sfix19_En18 
  input [18:0] Wgt_8_188, // sfix19_En18 
  input [18:0] Wgt_8_189, // sfix19_En18 
  input [18:0] Wgt_8_190, // sfix19_En18 
  input [18:0] Wgt_8_191, // sfix19_En18 
  input [18:0] Wgt_8_192, // sfix19_En18 
  input [18:0] Wgt_8_193, // sfix19_En18 
  input [18:0] Wgt_8_194, // sfix19_En18 
  input [18:0] Wgt_8_195, // sfix19_En18 
  input [18:0] Wgt_8_196, // sfix19_En18 
  input [18:0] Wgt_8_197, // sfix19_En18 
  input [18:0] Wgt_8_198, // sfix19_En18 
  input [18:0] Wgt_8_199, // sfix19_En18 
  input [18:0] Wgt_8_200, // sfix19_En18 
  input [18:0] Wgt_8_201, // sfix19_En18 
  input [18:0] Wgt_8_202, // sfix19_En18 
  input [18:0] Wgt_8_203, // sfix19_En18 
  input [18:0] Wgt_8_204, // sfix19_En18 
  input [18:0] Wgt_8_205, // sfix19_En18 
  input [18:0] Wgt_8_206, // sfix19_En18 
  input [18:0] Wgt_8_207, // sfix19_En18 
  input [18:0] Wgt_8_208, // sfix19_En18 
  input [18:0] Wgt_8_209, // sfix19_En18 
  input [18:0] Wgt_8_210, // sfix19_En18 
  input [18:0] Wgt_8_211, // sfix19_En18 
  input [18:0] Wgt_8_212, // sfix19_En18 
  input [18:0] Wgt_8_213, // sfix19_En18 
  input [18:0] Wgt_8_214, // sfix19_En18 
  input [18:0] Wgt_8_215, // sfix19_En18 
  input [18:0] Wgt_8_216, // sfix19_En18 
  input [18:0] Wgt_8_217, // sfix19_En18 
  input [18:0] Wgt_8_218, // sfix19_En18 
  input [18:0] Wgt_8_219, // sfix19_En18 
  input [18:0] Wgt_8_220, // sfix19_En18 
  input [18:0] Wgt_8_221, // sfix19_En18 
  input [18:0] Wgt_8_222, // sfix19_En18 
  input [18:0] Wgt_8_223, // sfix19_En18 
  input [18:0] Wgt_8_224, // sfix19_En18 
  input [18:0] Wgt_8_225, // sfix19_En18 
  input [18:0] Wgt_8_226, // sfix19_En18 
  input [18:0] Wgt_8_227, // sfix19_En18 
  input [18:0] Wgt_8_228, // sfix19_En18 
  input [18:0] Wgt_8_229, // sfix19_En18 
  input [18:0] Wgt_8_230, // sfix19_En18 
  input [18:0] Wgt_8_231, // sfix19_En18 
  input [18:0] Wgt_8_232, // sfix19_En18 
  input [18:0] Wgt_8_233, // sfix19_En18 
  input [18:0] Wgt_8_234, // sfix19_En18 
  input [18:0] Wgt_8_235, // sfix19_En18 
  input [18:0] Wgt_8_236, // sfix19_En18 
  input [18:0] Wgt_8_237, // sfix19_En18 
  input [18:0] Wgt_8_238, // sfix19_En18 
  input [18:0] Wgt_8_239, // sfix19_En18 
  input [18:0] Wgt_8_240, // sfix19_En18 
  input [18:0] Wgt_8_241, // sfix19_En18 
  input [18:0] Wgt_8_242, // sfix19_En18 
  input [18:0] Wgt_8_243, // sfix19_En18 
  input [18:0] Wgt_8_244, // sfix19_En18 
  input [18:0] Wgt_8_245, // sfix19_En18 
  input [18:0] Wgt_8_246, // sfix19_En18 
  input [18:0] Wgt_8_247, // sfix19_En18 
  input [18:0] Wgt_8_248, // sfix19_En18 
  input [18:0] Wgt_8_249, // sfix19_En18 
  input [18:0] Wgt_8_250, // sfix19_En18 
  input [18:0] Wgt_8_251, // sfix19_En18 
  input [18:0] Wgt_8_252, // sfix19_En18 
  input [18:0] Wgt_8_253, // sfix19_En18 
  input [18:0] Wgt_8_254, // sfix19_En18 
  input [18:0] Wgt_8_255, // sfix19_En18 
  input [18:0] Wgt_8_256, // sfix19_En18 
  input [18:0] Wgt_8_257, // sfix19_En18 
  input [18:0] Wgt_8_258, // sfix19_En18 
  input [18:0] Wgt_8_259, // sfix19_En18 
  input [18:0] Wgt_8_260, // sfix19_En18 
  input [18:0] Wgt_8_261, // sfix19_En18 
  input [18:0] Wgt_8_262, // sfix19_En18 
  input [18:0] Wgt_8_263, // sfix19_En18 
  input [18:0] Wgt_8_264, // sfix19_En18 
  input [18:0] Wgt_8_265, // sfix19_En18 
  input [18:0] Wgt_8_266, // sfix19_En18 
  input [18:0] Wgt_8_267, // sfix19_En18 
  input [18:0] Wgt_8_268, // sfix19_En18 
  input [18:0] Wgt_8_269, // sfix19_En18 
  input [18:0] Wgt_8_270, // sfix19_En18 
  input [18:0] Wgt_8_271, // sfix19_En18 
  input [18:0] Wgt_8_272, // sfix19_En18 
  input [18:0] Wgt_8_273, // sfix19_En18 
  input [18:0] Wgt_8_274, // sfix19_En18 
  input [18:0] Wgt_8_275, // sfix19_En18 
  input [18:0] Wgt_8_276, // sfix19_En18 
  input [18:0] Wgt_8_277, // sfix19_En18 
  input [18:0] Wgt_8_278, // sfix19_En18 
  input [18:0] Wgt_8_279, // sfix19_En18 
  input [18:0] Wgt_8_280, // sfix19_En18 
  input [18:0] Wgt_8_281, // sfix19_En18 
  input [18:0] Wgt_8_282, // sfix19_En18 
  input [18:0] Wgt_8_283, // sfix19_En18 
  input [18:0] Wgt_8_284, // sfix19_En18 
  input [18:0] Wgt_8_285, // sfix19_En18 
  input [18:0] Wgt_8_286, // sfix19_En18 
  input [18:0] Wgt_8_287, // sfix19_En18 
  input [18:0] Wgt_8_288, // sfix19_En18 
  input [18:0] Wgt_8_289, // sfix19_En18 
  input [18:0] Wgt_8_290, // sfix19_En18 
  input [18:0] Wgt_8_291, // sfix19_En18 
  input [18:0] Wgt_8_292, // sfix19_En18 
  input [18:0] Wgt_8_293, // sfix19_En18 
  input [18:0] Wgt_8_294, // sfix19_En18 
  input [18:0] Wgt_8_295, // sfix19_En18 
  input [18:0] Wgt_8_296, // sfix19_En18 
  input [18:0] Wgt_8_297, // sfix19_En18 
  input [18:0] Wgt_8_298, // sfix19_En18 
  input [18:0] Wgt_8_299, // sfix19_En18 
  input [18:0] Wgt_8_300, // sfix19_En18 
  input [18:0] Wgt_8_301, // sfix19_En18 
  input [18:0] Wgt_8_302, // sfix19_En18 
  input [18:0] Wgt_8_303, // sfix19_En18 
  input [18:0] Wgt_8_304, // sfix19_En18 
  input [18:0] Wgt_8_305, // sfix19_En18 
  input [18:0] Wgt_8_306, // sfix19_En18 
  input [18:0] Wgt_8_307, // sfix19_En18 
  input [18:0] Wgt_8_308, // sfix19_En18 
  input [18:0] Wgt_8_309, // sfix19_En18 
  input [18:0] Wgt_8_310, // sfix19_En18 
  input [18:0] Wgt_8_311, // sfix19_En18 
  input [18:0] Wgt_8_312, // sfix19_En18 
  input [18:0] Wgt_8_313, // sfix19_En18 
  input [18:0] Wgt_8_314, // sfix19_En18 
  input [18:0] Wgt_8_315, // sfix19_En18 
  input [18:0] Wgt_8_316, // sfix19_En18 
  input [18:0] Wgt_8_317, // sfix19_En18 
  input [18:0] Wgt_8_318, // sfix19_En18 
  input [18:0] Wgt_8_319, // sfix19_En18 
  input [18:0] Wgt_8_320, // sfix19_En18 
  input [18:0] Wgt_8_321, // sfix19_En18 
  input [18:0] Wgt_8_322, // sfix19_En18 
  input [18:0] Wgt_8_323, // sfix19_En18 
  input [18:0] Wgt_8_324, // sfix19_En18 
  input [18:0] Wgt_8_325, // sfix19_En18 
  input [18:0] Wgt_8_326, // sfix19_En18 
  input [18:0] Wgt_8_327, // sfix19_En18 
  input [18:0] Wgt_8_328, // sfix19_En18 
  input [18:0] Wgt_8_329, // sfix19_En18 
  input [18:0] Wgt_8_330, // sfix19_En18 
  input [18:0] Wgt_8_331, // sfix19_En18 
  input [18:0] Wgt_8_332, // sfix19_En18 
  input [18:0] Wgt_8_333, // sfix19_En18 
  input [18:0] Wgt_8_334, // sfix19_En18 
  input [18:0] Wgt_8_335, // sfix19_En18 
  input [18:0] Wgt_8_336, // sfix19_En18 
  input [18:0] Wgt_8_337, // sfix19_En18 
  input [18:0] Wgt_8_338, // sfix19_En18 
  input [18:0] Wgt_8_339, // sfix19_En18 
  input [18:0] Wgt_8_340, // sfix19_En18 
  input [18:0] Wgt_8_341, // sfix19_En18 
  input [18:0] Wgt_8_342, // sfix19_En18 
  input [18:0] Wgt_8_343, // sfix19_En18 
  input [18:0] Wgt_8_344, // sfix19_En18 
  input [18:0] Wgt_8_345, // sfix19_En18 
  input [18:0] Wgt_8_346, // sfix19_En18 
  input [18:0] Wgt_8_347, // sfix19_En18 
  input [18:0] Wgt_8_348, // sfix19_En18 
  input [18:0] Wgt_8_349, // sfix19_En18 
  input [18:0] Wgt_8_350, // sfix19_En18 
  input [18:0] Wgt_8_351, // sfix19_En18 
  input [18:0] Wgt_8_352, // sfix19_En18 
  input [18:0] Wgt_8_353, // sfix19_En18 
  input [18:0] Wgt_8_354, // sfix19_En18 
  input [18:0] Wgt_8_355, // sfix19_En18 
  input [18:0] Wgt_8_356, // sfix19_En18 
  input [18:0] Wgt_8_357, // sfix19_En18 
  input [18:0] Wgt_8_358, // sfix19_En18 
  input [18:0] Wgt_8_359, // sfix19_En18 
  input [18:0] Wgt_8_360, // sfix19_En18 
  input [18:0] Wgt_8_361, // sfix19_En18 
  input [18:0] Wgt_8_362, // sfix19_En18 
  input [18:0] Wgt_8_363, // sfix19_En18 
  input [18:0] Wgt_8_364, // sfix19_En18 
  input [18:0] Wgt_8_365, // sfix19_En18 
  input [18:0] Wgt_8_366, // sfix19_En18 
  input [18:0] Wgt_8_367, // sfix19_En18 
  input [18:0] Wgt_8_368, // sfix19_En18 
  input [18:0] Wgt_8_369, // sfix19_En18 
  input [18:0] Wgt_8_370, // sfix19_En18 
  input [18:0] Wgt_8_371, // sfix19_En18 
  input [18:0] Wgt_8_372, // sfix19_En18 
  input [18:0] Wgt_8_373, // sfix19_En18 
  input [18:0] Wgt_8_374, // sfix19_En18 
  input [18:0] Wgt_8_375, // sfix19_En18 
  input [18:0] Wgt_8_376, // sfix19_En18 
  input [18:0] Wgt_8_377, // sfix19_En18 
  input [18:0] Wgt_8_378, // sfix19_En18 
  input [18:0] Wgt_8_379, // sfix19_En18 
  input [18:0] Wgt_8_380, // sfix19_En18 
  input [18:0] Wgt_8_381, // sfix19_En18 
  input [18:0] Wgt_8_382, // sfix19_En18 
  input [18:0] Wgt_8_383, // sfix19_En18 
  input [18:0] Wgt_8_384, // sfix19_En18 
  input [18:0] Wgt_8_385, // sfix19_En18 
  input [18:0] Wgt_8_386, // sfix19_En18 
  input [18:0] Wgt_8_387, // sfix19_En18 
  input [18:0] Wgt_8_388, // sfix19_En18 
  input [18:0] Wgt_8_389, // sfix19_En18 
  input [18:0] Wgt_8_390, // sfix19_En18 
  input [18:0] Wgt_8_391, // sfix19_En18 
  input [18:0] Wgt_8_392, // sfix19_En18 
  input [18:0] Wgt_8_393, // sfix19_En18 
  input [18:0] Wgt_8_394, // sfix19_En18 
  input [18:0] Wgt_8_395, // sfix19_En18 
  input [18:0] Wgt_8_396, // sfix19_En18 
  input [18:0] Wgt_8_397, // sfix19_En18 
  input [18:0] Wgt_8_398, // sfix19_En18 
  input [18:0] Wgt_8_399, // sfix19_En18 
  input [18:0] Wgt_8_400, // sfix19_En18 
  input [18:0] Wgt_8_401, // sfix19_En18 
  input [18:0] Wgt_8_402, // sfix19_En18 
  input [18:0] Wgt_8_403, // sfix19_En18 
  input [18:0] Wgt_8_404, // sfix19_En18 
  input [18:0] Wgt_8_405, // sfix19_En18 
  input [18:0] Wgt_8_406, // sfix19_En18 
  input [18:0] Wgt_8_407, // sfix19_En18 
  input [18:0] Wgt_8_408, // sfix19_En18 
  input [18:0] Wgt_8_409, // sfix19_En18 
  input [18:0] Wgt_8_410, // sfix19_En18 
  input [18:0] Wgt_8_411, // sfix19_En18 
  input [18:0] Wgt_8_412, // sfix19_En18 
  input [18:0] Wgt_8_413, // sfix19_En18 
  input [18:0] Wgt_8_414, // sfix19_En18 
  input [18:0] Wgt_8_415, // sfix19_En18 
  input [18:0] Wgt_8_416, // sfix19_En18 
  input [18:0] Wgt_8_417, // sfix19_En18 
  input [18:0] Wgt_8_418, // sfix19_En18 
  input [18:0] Wgt_8_419, // sfix19_En18 
  input [18:0] Wgt_8_420, // sfix19_En18 
  input [18:0] Wgt_8_421, // sfix19_En18 
  input [18:0] Wgt_8_422, // sfix19_En18 
  input [18:0] Wgt_8_423, // sfix19_En18 
  input [18:0] Wgt_8_424, // sfix19_En18 
  input [18:0] Wgt_8_425, // sfix19_En18 
  input [18:0] Wgt_8_426, // sfix19_En18 
  input [18:0] Wgt_8_427, // sfix19_En18 
  input [18:0] Wgt_8_428, // sfix19_En18 
  input [18:0] Wgt_8_429, // sfix19_En18 
  input [18:0] Wgt_8_430, // sfix19_En18 
  input [18:0] Wgt_8_431, // sfix19_En18 
  input [18:0] Wgt_8_432, // sfix19_En18 
  input [18:0] Wgt_8_433, // sfix19_En18 
  input [18:0] Wgt_8_434, // sfix19_En18 
  input [18:0] Wgt_8_435, // sfix19_En18 
  input [18:0] Wgt_8_436, // sfix19_En18 
  input [18:0] Wgt_8_437, // sfix19_En18 
  input [18:0] Wgt_8_438, // sfix19_En18 
  input [18:0] Wgt_8_439, // sfix19_En18 
  input [18:0] Wgt_8_440, // sfix19_En18 
  input [18:0] Wgt_8_441, // sfix19_En18 
  input [18:0] Wgt_8_442, // sfix19_En18 
  input [18:0] Wgt_8_443, // sfix19_En18 
  input [18:0] Wgt_8_444, // sfix19_En18 
  input [18:0] Wgt_8_445, // sfix19_En18 
  input [18:0] Wgt_8_446, // sfix19_En18 
  input [18:0] Wgt_8_447, // sfix19_En18 
  input [18:0] Wgt_8_448, // sfix19_En18 
  input [18:0] Wgt_8_449, // sfix19_En18 
  input [18:0] Wgt_8_450, // sfix19_En18 
  input [18:0] Wgt_8_451, // sfix19_En18 
  input [18:0] Wgt_8_452, // sfix19_En18 
  input [18:0] Wgt_8_453, // sfix19_En18 
  input [18:0] Wgt_8_454, // sfix19_En18 
  input [18:0] Wgt_8_455, // sfix19_En18 
  input [18:0] Wgt_8_456, // sfix19_En18 
  input [18:0] Wgt_8_457, // sfix19_En18 
  input [18:0] Wgt_8_458, // sfix19_En18 
  input [18:0] Wgt_8_459, // sfix19_En18 
  input [18:0] Wgt_8_460, // sfix19_En18 
  input [18:0] Wgt_8_461, // sfix19_En18 
  input [18:0] Wgt_8_462, // sfix19_En18 
  input [18:0] Wgt_8_463, // sfix19_En18 
  input [18:0] Wgt_8_464, // sfix19_En18 
  input [18:0] Wgt_8_465, // sfix19_En18 
  input [18:0] Wgt_8_466, // sfix19_En18 
  input [18:0] Wgt_8_467, // sfix19_En18 
  input [18:0] Wgt_8_468, // sfix19_En18 
  input [18:0] Wgt_8_469, // sfix19_En18 
  input [18:0] Wgt_8_470, // sfix19_En18 
  input [18:0] Wgt_8_471, // sfix19_En18 
  input [18:0] Wgt_8_472, // sfix19_En18 
  input [18:0] Wgt_8_473, // sfix19_En18 
  input [18:0] Wgt_8_474, // sfix19_En18 
  input [18:0] Wgt_8_475, // sfix19_En18 
  input [18:0] Wgt_8_476, // sfix19_En18 
  input [18:0] Wgt_8_477, // sfix19_En18 
  input [18:0] Wgt_8_478, // sfix19_En18 
  input [18:0] Wgt_8_479, // sfix19_En18 
  input [18:0] Wgt_8_480, // sfix19_En18 
  input [18:0] Wgt_8_481, // sfix19_En18 
  input [18:0] Wgt_8_482, // sfix19_En18 
  input [18:0] Wgt_8_483, // sfix19_En18 
  input [18:0] Wgt_8_484, // sfix19_En18 
  input [18:0] Wgt_8_485, // sfix19_En18 
  input [18:0] Wgt_8_486, // sfix19_En18 
  input [18:0] Wgt_8_487, // sfix19_En18 
  input [18:0] Wgt_8_488, // sfix19_En18 
  input [18:0] Wgt_8_489, // sfix19_En18 
  input [18:0] Wgt_8_490, // sfix19_En18 
  input [18:0] Wgt_8_491, // sfix19_En18 
  input [18:0] Wgt_8_492, // sfix19_En18 
  input [18:0] Wgt_8_493, // sfix19_En18 
  input [18:0] Wgt_8_494, // sfix19_En18 
  input [18:0] Wgt_8_495, // sfix19_En18 
  input [18:0] Wgt_8_496, // sfix19_En18 
  input [18:0] Wgt_8_497, // sfix19_En18 
  input [18:0] Wgt_8_498, // sfix19_En18 
  input [18:0] Wgt_8_499, // sfix19_En18 
  input [18:0] Wgt_8_500, // sfix19_En18 
  input [18:0] Wgt_8_501, // sfix19_En18 
  input [18:0] Wgt_8_502, // sfix19_En18 
  input [18:0] Wgt_8_503, // sfix19_En18 
  input [18:0] Wgt_8_504, // sfix19_En18 
  input [18:0] Wgt_8_505, // sfix19_En18 
  input [18:0] Wgt_8_506, // sfix19_En18 
  input [18:0] Wgt_8_507, // sfix19_En18 
  input [18:0] Wgt_8_508, // sfix19_En18 
  input [18:0] Wgt_8_509, // sfix19_En18 
  input [18:0] Wgt_8_510, // sfix19_En18 
  input [18:0] Wgt_8_511, // sfix19_En18 
  input [18:0] Wgt_8_512, // sfix19_En18 
  input [18:0] Wgt_8_513, // sfix19_En18 
  input [18:0] Wgt_8_514, // sfix19_En18 
  input [18:0] Wgt_8_515, // sfix19_En18 
  input [18:0] Wgt_8_516, // sfix19_En18 
  input [18:0] Wgt_8_517, // sfix19_En18 
  input [18:0] Wgt_8_518, // sfix19_En18 
  input [18:0] Wgt_8_519, // sfix19_En18 
  input [18:0] Wgt_8_520, // sfix19_En18 
  input [18:0] Wgt_8_521, // sfix19_En18 
  input [18:0] Wgt_8_522, // sfix19_En18 
  input [18:0] Wgt_8_523, // sfix19_En18 
  input [18:0] Wgt_8_524, // sfix19_En18 
  input [18:0] Wgt_8_525, // sfix19_En18 
  input [18:0] Wgt_8_526, // sfix19_En18 
  input [18:0] Wgt_8_527, // sfix19_En18 
  input [18:0] Wgt_8_528, // sfix19_En18 
  input [18:0] Wgt_8_529, // sfix19_En18 
  input [18:0] Wgt_8_530, // sfix19_En18 
  input [18:0] Wgt_8_531, // sfix19_En18 
  input [18:0] Wgt_8_532, // sfix19_En18 
  input [18:0] Wgt_8_533, // sfix19_En18 
  input [18:0] Wgt_8_534, // sfix19_En18 
  input [18:0] Wgt_8_535, // sfix19_En18 
  input [18:0] Wgt_8_536, // sfix19_En18 
  input [18:0] Wgt_8_537, // sfix19_En18 
  input [18:0] Wgt_8_538, // sfix19_En18 
  input [18:0] Wgt_8_539, // sfix19_En18 
  input [18:0] Wgt_8_540, // sfix19_En18 
  input [18:0] Wgt_8_541, // sfix19_En18 
  input [18:0] Wgt_8_542, // sfix19_En18 
  input [18:0] Wgt_8_543, // sfix19_En18 
  input [18:0] Wgt_8_544, // sfix19_En18 
  input [18:0] Wgt_8_545, // sfix19_En18 
  input [18:0] Wgt_8_546, // sfix19_En18 
  input [18:0] Wgt_8_547, // sfix19_En18 
  input [18:0] Wgt_8_548, // sfix19_En18 
  input [18:0] Wgt_8_549, // sfix19_En18 
  input [18:0] Wgt_8_550, // sfix19_En18 
  input [18:0] Wgt_8_551, // sfix19_En18 
  input [18:0] Wgt_8_552, // sfix19_En18 
  input [18:0] Wgt_8_553, // sfix19_En18 
  input [18:0] Wgt_8_554, // sfix19_En18 
  input [18:0] Wgt_8_555, // sfix19_En18 
  input [18:0] Wgt_8_556, // sfix19_En18 
  input [18:0] Wgt_8_557, // sfix19_En18 
  input [18:0] Wgt_8_558, // sfix19_En18 
  input [18:0] Wgt_8_559, // sfix19_En18 
  input [18:0] Wgt_8_560, // sfix19_En18 
  input [18:0] Wgt_8_561, // sfix19_En18 
  input [18:0] Wgt_8_562, // sfix19_En18 
  input [18:0] Wgt_8_563, // sfix19_En18 
  input [18:0] Wgt_8_564, // sfix19_En18 
  input [18:0] Wgt_8_565, // sfix19_En18 
  input [18:0] Wgt_8_566, // sfix19_En18 
  input [18:0] Wgt_8_567, // sfix19_En18 
  input [18:0] Wgt_8_568, // sfix19_En18 
  input [18:0] Wgt_8_569, // sfix19_En18 
  input [18:0] Wgt_8_570, // sfix19_En18 
  input [18:0] Wgt_8_571, // sfix19_En18 
  input [18:0] Wgt_8_572, // sfix19_En18 
  input [18:0] Wgt_8_573, // sfix19_En18 
  input [18:0] Wgt_8_574, // sfix19_En18 
  input [18:0] Wgt_8_575, // sfix19_En18 
  input [18:0] Wgt_8_576, // sfix19_En18 
  input [18:0] Wgt_8_577, // sfix19_En18 
  input [18:0] Wgt_8_578, // sfix19_En18 
  input [18:0] Wgt_8_579, // sfix19_En18 
  input [18:0] Wgt_8_580, // sfix19_En18 
  input [18:0] Wgt_8_581, // sfix19_En18 
  input [18:0] Wgt_8_582, // sfix19_En18 
  input [18:0] Wgt_8_583, // sfix19_En18 
  input [18:0] Wgt_8_584, // sfix19_En18 
  input [18:0] Wgt_8_585, // sfix19_En18 
  input [18:0] Wgt_8_586, // sfix19_En18 
  input [18:0] Wgt_8_587, // sfix19_En18 
  input [18:0] Wgt_8_588, // sfix19_En18 
  input [18:0] Wgt_8_589, // sfix19_En18 
  input [18:0] Wgt_8_590, // sfix19_En18 
  input [18:0] Wgt_8_591, // sfix19_En18 
  input [18:0] Wgt_8_592, // sfix19_En18 
  input [18:0] Wgt_8_593, // sfix19_En18 
  input [18:0] Wgt_8_594, // sfix19_En18 
  input [18:0] Wgt_8_595, // sfix19_En18 
  input [18:0] Wgt_8_596, // sfix19_En18 
  input [18:0] Wgt_8_597, // sfix19_En18 
  input [18:0] Wgt_8_598, // sfix19_En18 
  input [18:0] Wgt_8_599, // sfix19_En18 
  input [18:0] Wgt_8_600, // sfix19_En18 
  input [18:0] Wgt_8_601, // sfix19_En18 
  input [18:0] Wgt_8_602, // sfix19_En18 
  input [18:0] Wgt_8_603, // sfix19_En18 
  input [18:0] Wgt_8_604, // sfix19_En18 
  input [18:0] Wgt_8_605, // sfix19_En18 
  input [18:0] Wgt_8_606, // sfix19_En18 
  input [18:0] Wgt_8_607, // sfix19_En18 
  input [18:0] Wgt_8_608, // sfix19_En18 
  input [18:0] Wgt_8_609, // sfix19_En18 
  input [18:0] Wgt_8_610, // sfix19_En18 
  input [18:0] Wgt_8_611, // sfix19_En18 
  input [18:0] Wgt_8_612, // sfix19_En18 
  input [18:0] Wgt_8_613, // sfix19_En18 
  input [18:0] Wgt_8_614, // sfix19_En18 
  input [18:0] Wgt_8_615, // sfix19_En18 
  input [18:0] Wgt_8_616, // sfix19_En18 
  input [18:0] Wgt_8_617, // sfix19_En18 
  input [18:0] Wgt_8_618, // sfix19_En18 
  input [18:0] Wgt_8_619, // sfix19_En18 
  input [18:0] Wgt_8_620, // sfix19_En18 
  input [18:0] Wgt_8_621, // sfix19_En18 
  input [18:0] Wgt_8_622, // sfix19_En18 
  input [18:0] Wgt_8_623, // sfix19_En18 
  input [18:0] Wgt_8_624, // sfix19_En18 
  input [18:0] Wgt_8_625, // sfix19_En18 
  input [18:0] Wgt_8_626, // sfix19_En18 
  input [18:0] Wgt_8_627, // sfix19_En18 
  input [18:0] Wgt_8_628, // sfix19_En18 
  input [18:0] Wgt_8_629, // sfix19_En18 
  input [18:0] Wgt_8_630, // sfix19_En18 
  input [18:0] Wgt_8_631, // sfix19_En18 
  input [18:0] Wgt_8_632, // sfix19_En18 
  input [18:0] Wgt_8_633, // sfix19_En18 
  input [18:0] Wgt_8_634, // sfix19_En18 
  input [18:0] Wgt_8_635, // sfix19_En18 
  input [18:0] Wgt_8_636, // sfix19_En18 
  input [18:0] Wgt_8_637, // sfix19_En18 
  input [18:0] Wgt_8_638, // sfix19_En18 
  input [18:0] Wgt_8_639, // sfix19_En18 
  input [18:0] Wgt_8_640, // sfix19_En18 
  input [18:0] Wgt_8_641, // sfix19_En18 
  input [18:0] Wgt_8_642, // sfix19_En18 
  input [18:0] Wgt_8_643, // sfix19_En18 
  input [18:0] Wgt_8_644, // sfix19_En18 
  input [18:0] Wgt_8_645, // sfix19_En18 
  input [18:0] Wgt_8_646, // sfix19_En18 
  input [18:0] Wgt_8_647, // sfix19_En18 
  input [18:0] Wgt_8_648, // sfix19_En18 
  input [18:0] Wgt_8_649, // sfix19_En18 
  input [18:0] Wgt_8_650, // sfix19_En18 
  input [18:0] Wgt_8_651, // sfix19_En18 
  input [18:0] Wgt_8_652, // sfix19_En18 
  input [18:0] Wgt_8_653, // sfix19_En18 
  input [18:0] Wgt_8_654, // sfix19_En18 
  input [18:0] Wgt_8_655, // sfix19_En18 
  input [18:0] Wgt_8_656, // sfix19_En18 
  input [18:0] Wgt_8_657, // sfix19_En18 
  input [18:0] Wgt_8_658, // sfix19_En18 
  input [18:0] Wgt_8_659, // sfix19_En18 
  input [18:0] Wgt_8_660, // sfix19_En18 
  input [18:0] Wgt_8_661, // sfix19_En18 
  input [18:0] Wgt_8_662, // sfix19_En18 
  input [18:0] Wgt_8_663, // sfix19_En18 
  input [18:0] Wgt_8_664, // sfix19_En18 
  input [18:0] Wgt_8_665, // sfix19_En18 
  input [18:0] Wgt_8_666, // sfix19_En18 
  input [18:0] Wgt_8_667, // sfix19_En18 
  input [18:0] Wgt_8_668, // sfix19_En18 
  input [18:0] Wgt_8_669, // sfix19_En18 
  input [18:0] Wgt_8_670, // sfix19_En18 
  input [18:0] Wgt_8_671, // sfix19_En18 
  input [18:0] Wgt_8_672, // sfix19_En18 
  input [18:0] Wgt_8_673, // sfix19_En18 
  input [18:0] Wgt_8_674, // sfix19_En18 
  input [18:0] Wgt_8_675, // sfix19_En18 
  input [18:0] Wgt_8_676, // sfix19_En18 
  input [18:0] Wgt_8_677, // sfix19_En18 
  input [18:0] Wgt_8_678, // sfix19_En18 
  input [18:0] Wgt_8_679, // sfix19_En18 
  input [18:0] Wgt_8_680, // sfix19_En18 
  input [18:0] Wgt_8_681, // sfix19_En18 
  input [18:0] Wgt_8_682, // sfix19_En18 
  input [18:0] Wgt_8_683, // sfix19_En18 
  input [18:0] Wgt_8_684, // sfix19_En18 
  input [18:0] Wgt_8_685, // sfix19_En18 
  input [18:0] Wgt_8_686, // sfix19_En18 
  input [18:0] Wgt_8_687, // sfix19_En18 
  input [18:0] Wgt_8_688, // sfix19_En18 
  input [18:0] Wgt_8_689, // sfix19_En18 
  input [18:0] Wgt_8_690, // sfix19_En18 
  input [18:0] Wgt_8_691, // sfix19_En18 
  input [18:0] Wgt_8_692, // sfix19_En18 
  input [18:0] Wgt_8_693, // sfix19_En18 
  input [18:0] Wgt_8_694, // sfix19_En18 
  input [18:0] Wgt_8_695, // sfix19_En18 
  input [18:0] Wgt_8_696, // sfix19_En18 
  input [18:0] Wgt_8_697, // sfix19_En18 
  input [18:0] Wgt_8_698, // sfix19_En18 
  input [18:0] Wgt_8_699, // sfix19_En18 
  input [18:0] Wgt_8_700, // sfix19_En18 
  input [18:0] Wgt_8_701, // sfix19_En18 
  input [18:0] Wgt_8_702, // sfix19_En18 
  input [18:0] Wgt_8_703, // sfix19_En18 
  input [18:0] Wgt_8_704, // sfix19_En18 
  input [18:0] Wgt_8_705, // sfix19_En18 
  input [18:0] Wgt_8_706, // sfix19_En18 
  input [18:0] Wgt_8_707, // sfix19_En18 
  input [18:0] Wgt_8_708, // sfix19_En18 
  input [18:0] Wgt_8_709, // sfix19_En18 
  input [18:0] Wgt_8_710, // sfix19_En18 
  input [18:0] Wgt_8_711, // sfix19_En18 
  input [18:0] Wgt_8_712, // sfix19_En18 
  input [18:0] Wgt_8_713, // sfix19_En18 
  input [18:0] Wgt_8_714, // sfix19_En18 
  input [18:0] Wgt_8_715, // sfix19_En18 
  input [18:0] Wgt_8_716, // sfix19_En18 
  input [18:0] Wgt_8_717, // sfix19_En18 
  input [18:0] Wgt_8_718, // sfix19_En18 
  input [18:0] Wgt_8_719, // sfix19_En18 
  input [18:0] Wgt_8_720, // sfix19_En18 
  input [18:0] Wgt_8_721, // sfix19_En18 
  input [18:0] Wgt_8_722, // sfix19_En18 
  input [18:0] Wgt_8_723, // sfix19_En18 
  input [18:0] Wgt_8_724, // sfix19_En18 
  input [18:0] Wgt_8_725, // sfix19_En18 
  input [18:0] Wgt_8_726, // sfix19_En18 
  input [18:0] Wgt_8_727, // sfix19_En18 
  input [18:0] Wgt_8_728, // sfix19_En18 
  input [18:0] Wgt_8_729, // sfix19_En18 
  input [18:0] Wgt_8_730, // sfix19_En18 
  input [18:0] Wgt_8_731, // sfix19_En18 
  input [18:0] Wgt_8_732, // sfix19_En18 
  input [18:0] Wgt_8_733, // sfix19_En18 
  input [18:0] Wgt_8_734, // sfix19_En18 
  input [18:0] Wgt_8_735, // sfix19_En18 
  input [18:0] Wgt_8_736, // sfix19_En18 
  input [18:0] Wgt_8_737, // sfix19_En18 
  input [18:0] Wgt_8_738, // sfix19_En18 
  input [18:0] Wgt_8_739, // sfix19_En18 
  input [18:0] Wgt_8_740, // sfix19_En18 
  input [18:0] Wgt_8_741, // sfix19_En18 
  input [18:0] Wgt_8_742, // sfix19_En18 
  input [18:0] Wgt_8_743, // sfix19_En18 
  input [18:0] Wgt_8_744, // sfix19_En18 
  input [18:0] Wgt_8_745, // sfix19_En18 
  input [18:0] Wgt_8_746, // sfix19_En18 
  input [18:0] Wgt_8_747, // sfix19_En18 
  input [18:0] Wgt_8_748, // sfix19_En18 
  input [18:0] Wgt_8_749, // sfix19_En18 
  input [18:0] Wgt_8_750, // sfix19_En18 
  input [18:0] Wgt_8_751, // sfix19_En18 
  input [18:0] Wgt_8_752, // sfix19_En18 
  input [18:0] Wgt_8_753, // sfix19_En18 
  input [18:0] Wgt_8_754, // sfix19_En18 
  input [18:0] Wgt_8_755, // sfix19_En18 
  input [18:0] Wgt_8_756, // sfix19_En18 
  input [18:0] Wgt_8_757, // sfix19_En18 
  input [18:0] Wgt_8_758, // sfix19_En18 
  input [18:0] Wgt_8_759, // sfix19_En18 
  input [18:0] Wgt_8_760, // sfix19_En18 
  input [18:0] Wgt_8_761, // sfix19_En18 
  input [18:0] Wgt_8_762, // sfix19_En18 
  input [18:0] Wgt_8_763, // sfix19_En18 
  input [18:0] Wgt_8_764, // sfix19_En18 
  input [18:0] Wgt_8_765, // sfix19_En18 
  input [18:0] Wgt_8_766, // sfix19_En18 
  input [18:0] Wgt_8_767, // sfix19_En18 
  input [18:0] Wgt_8_768, // sfix19_En18 
  input [18:0] Wgt_8_769, // sfix19_En18 
  input [18:0] Wgt_8_770, // sfix19_En18 
  input [18:0] Wgt_8_771, // sfix19_En18 
  input [18:0] Wgt_8_772, // sfix19_En18 
  input [18:0] Wgt_8_773, // sfix19_En18 
  input [18:0] Wgt_8_774, // sfix19_En18 
  input [18:0] Wgt_8_775, // sfix19_En18 
  input [18:0] Wgt_8_776, // sfix19_En18 
  input [18:0] Wgt_8_777, // sfix19_En18 
  input [18:0] Wgt_8_778, // sfix19_En18 
  input [18:0] Wgt_8_779, // sfix19_En18 
  input [18:0] Wgt_8_780, // sfix19_En18 
  input [18:0] Wgt_8_781, // sfix19_En18 
  input [18:0] Wgt_8_782, // sfix19_En18 
  input [18:0] Wgt_8_783, // sfix19_En18 
  input [18:0] Wgt_8_784, // sfix19_En18 
  input [18:0] Wgt_9_0, // sfix19_En18 
  input [18:0] Wgt_9_1, // sfix19_En18 
  input [18:0] Wgt_9_2, // sfix19_En18 
  input [18:0] Wgt_9_3, // sfix19_En18 
  input [18:0] Wgt_9_4, // sfix19_En18 
  input [18:0] Wgt_9_5, // sfix19_En18 
  input [18:0] Wgt_9_6, // sfix19_En18 
  input [18:0] Wgt_9_7, // sfix19_En18 
  input [18:0] Wgt_9_8, // sfix19_En18 
  input [18:0] Wgt_9_9, // sfix19_En18 
  input [18:0] Wgt_9_10, // sfix19_En18 
  input [18:0] Wgt_9_11, // sfix19_En18 
  input [18:0] Wgt_9_12, // sfix19_En18 
  input [18:0] Wgt_9_13, // sfix19_En18 
  input [18:0] Wgt_9_14, // sfix19_En18 
  input [18:0] Wgt_9_15, // sfix19_En18 
  input [18:0] Wgt_9_16, // sfix19_En18 
  input [18:0] Wgt_9_17, // sfix19_En18 
  input [18:0] Wgt_9_18, // sfix19_En18 
  input [18:0] Wgt_9_19, // sfix19_En18 
  input [18:0] Wgt_9_20, // sfix19_En18 
  input [18:0] Wgt_9_21, // sfix19_En18 
  input [18:0] Wgt_9_22, // sfix19_En18 
  input [18:0] Wgt_9_23, // sfix19_En18 
  input [18:0] Wgt_9_24, // sfix19_En18 
  input [18:0] Wgt_9_25, // sfix19_En18 
  input [18:0] Wgt_9_26, // sfix19_En18 
  input [18:0] Wgt_9_27, // sfix19_En18 
  input [18:0] Wgt_9_28, // sfix19_En18 
  input [18:0] Wgt_9_29, // sfix19_En18 
  input [18:0] Wgt_9_30, // sfix19_En18 
  input [18:0] Wgt_9_31, // sfix19_En18 
  input [18:0] Wgt_9_32, // sfix19_En18 
  input [18:0] Wgt_9_33, // sfix19_En18 
  input [18:0] Wgt_9_34, // sfix19_En18 
  input [18:0] Wgt_9_35, // sfix19_En18 
  input [18:0] Wgt_9_36, // sfix19_En18 
  input [18:0] Wgt_9_37, // sfix19_En18 
  input [18:0] Wgt_9_38, // sfix19_En18 
  input [18:0] Wgt_9_39, // sfix19_En18 
  input [18:0] Wgt_9_40, // sfix19_En18 
  input [18:0] Wgt_9_41, // sfix19_En18 
  input [18:0] Wgt_9_42, // sfix19_En18 
  input [18:0] Wgt_9_43, // sfix19_En18 
  input [18:0] Wgt_9_44, // sfix19_En18 
  input [18:0] Wgt_9_45, // sfix19_En18 
  input [18:0] Wgt_9_46, // sfix19_En18 
  input [18:0] Wgt_9_47, // sfix19_En18 
  input [18:0] Wgt_9_48, // sfix19_En18 
  input [18:0] Wgt_9_49, // sfix19_En18 
  input [18:0] Wgt_9_50, // sfix19_En18 
  input [18:0] Wgt_9_51, // sfix19_En18 
  input [18:0] Wgt_9_52, // sfix19_En18 
  input [18:0] Wgt_9_53, // sfix19_En18 
  input [18:0] Wgt_9_54, // sfix19_En18 
  input [18:0] Wgt_9_55, // sfix19_En18 
  input [18:0] Wgt_9_56, // sfix19_En18 
  input [18:0] Wgt_9_57, // sfix19_En18 
  input [18:0] Wgt_9_58, // sfix19_En18 
  input [18:0] Wgt_9_59, // sfix19_En18 
  input [18:0] Wgt_9_60, // sfix19_En18 
  input [18:0] Wgt_9_61, // sfix19_En18 
  input [18:0] Wgt_9_62, // sfix19_En18 
  input [18:0] Wgt_9_63, // sfix19_En18 
  input [18:0] Wgt_9_64, // sfix19_En18 
  input [18:0] Wgt_9_65, // sfix19_En18 
  input [18:0] Wgt_9_66, // sfix19_En18 
  input [18:0] Wgt_9_67, // sfix19_En18 
  input [18:0] Wgt_9_68, // sfix19_En18 
  input [18:0] Wgt_9_69, // sfix19_En18 
  input [18:0] Wgt_9_70, // sfix19_En18 
  input [18:0] Wgt_9_71, // sfix19_En18 
  input [18:0] Wgt_9_72, // sfix19_En18 
  input [18:0] Wgt_9_73, // sfix19_En18 
  input [18:0] Wgt_9_74, // sfix19_En18 
  input [18:0] Wgt_9_75, // sfix19_En18 
  input [18:0] Wgt_9_76, // sfix19_En18 
  input [18:0] Wgt_9_77, // sfix19_En18 
  input [18:0] Wgt_9_78, // sfix19_En18 
  input [18:0] Wgt_9_79, // sfix19_En18 
  input [18:0] Wgt_9_80, // sfix19_En18 
  input [18:0] Wgt_9_81, // sfix19_En18 
  input [18:0] Wgt_9_82, // sfix19_En18 
  input [18:0] Wgt_9_83, // sfix19_En18 
  input [18:0] Wgt_9_84, // sfix19_En18 
  input [18:0] Wgt_9_85, // sfix19_En18 
  input [18:0] Wgt_9_86, // sfix19_En18 
  input [18:0] Wgt_9_87, // sfix19_En18 
  input [18:0] Wgt_9_88, // sfix19_En18 
  input [18:0] Wgt_9_89, // sfix19_En18 
  input [18:0] Wgt_9_90, // sfix19_En18 
  input [18:0] Wgt_9_91, // sfix19_En18 
  input [18:0] Wgt_9_92, // sfix19_En18 
  input [18:0] Wgt_9_93, // sfix19_En18 
  input [18:0] Wgt_9_94, // sfix19_En18 
  input [18:0] Wgt_9_95, // sfix19_En18 
  input [18:0] Wgt_9_96, // sfix19_En18 
  input [18:0] Wgt_9_97, // sfix19_En18 
  input [18:0] Wgt_9_98, // sfix19_En18 
  input [18:0] Wgt_9_99, // sfix19_En18 
  input [18:0] Wgt_9_100, // sfix19_En18 
  input [18:0] Wgt_9_101, // sfix19_En18 
  input [18:0] Wgt_9_102, // sfix19_En18 
  input [18:0] Wgt_9_103, // sfix19_En18 
  input [18:0] Wgt_9_104, // sfix19_En18 
  input [18:0] Wgt_9_105, // sfix19_En18 
  input [18:0] Wgt_9_106, // sfix19_En18 
  input [18:0] Wgt_9_107, // sfix19_En18 
  input [18:0] Wgt_9_108, // sfix19_En18 
  input [18:0] Wgt_9_109, // sfix19_En18 
  input [18:0] Wgt_9_110, // sfix19_En18 
  input [18:0] Wgt_9_111, // sfix19_En18 
  input [18:0] Wgt_9_112, // sfix19_En18 
  input [18:0] Wgt_9_113, // sfix19_En18 
  input [18:0] Wgt_9_114, // sfix19_En18 
  input [18:0] Wgt_9_115, // sfix19_En18 
  input [18:0] Wgt_9_116, // sfix19_En18 
  input [18:0] Wgt_9_117, // sfix19_En18 
  input [18:0] Wgt_9_118, // sfix19_En18 
  input [18:0] Wgt_9_119, // sfix19_En18 
  input [18:0] Wgt_9_120, // sfix19_En18 
  input [18:0] Wgt_9_121, // sfix19_En18 
  input [18:0] Wgt_9_122, // sfix19_En18 
  input [18:0] Wgt_9_123, // sfix19_En18 
  input [18:0] Wgt_9_124, // sfix19_En18 
  input [18:0] Wgt_9_125, // sfix19_En18 
  input [18:0] Wgt_9_126, // sfix19_En18 
  input [18:0] Wgt_9_127, // sfix19_En18 
  input [18:0] Wgt_9_128, // sfix19_En18 
  input [18:0] Wgt_9_129, // sfix19_En18 
  input [18:0] Wgt_9_130, // sfix19_En18 
  input [18:0] Wgt_9_131, // sfix19_En18 
  input [18:0] Wgt_9_132, // sfix19_En18 
  input [18:0] Wgt_9_133, // sfix19_En18 
  input [18:0] Wgt_9_134, // sfix19_En18 
  input [18:0] Wgt_9_135, // sfix19_En18 
  input [18:0] Wgt_9_136, // sfix19_En18 
  input [18:0] Wgt_9_137, // sfix19_En18 
  input [18:0] Wgt_9_138, // sfix19_En18 
  input [18:0] Wgt_9_139, // sfix19_En18 
  input [18:0] Wgt_9_140, // sfix19_En18 
  input [18:0] Wgt_9_141, // sfix19_En18 
  input [18:0] Wgt_9_142, // sfix19_En18 
  input [18:0] Wgt_9_143, // sfix19_En18 
  input [18:0] Wgt_9_144, // sfix19_En18 
  input [18:0] Wgt_9_145, // sfix19_En18 
  input [18:0] Wgt_9_146, // sfix19_En18 
  input [18:0] Wgt_9_147, // sfix19_En18 
  input [18:0] Wgt_9_148, // sfix19_En18 
  input [18:0] Wgt_9_149, // sfix19_En18 
  input [18:0] Wgt_9_150, // sfix19_En18 
  input [18:0] Wgt_9_151, // sfix19_En18 
  input [18:0] Wgt_9_152, // sfix19_En18 
  input [18:0] Wgt_9_153, // sfix19_En18 
  input [18:0] Wgt_9_154, // sfix19_En18 
  input [18:0] Wgt_9_155, // sfix19_En18 
  input [18:0] Wgt_9_156, // sfix19_En18 
  input [18:0] Wgt_9_157, // sfix19_En18 
  input [18:0] Wgt_9_158, // sfix19_En18 
  input [18:0] Wgt_9_159, // sfix19_En18 
  input [18:0] Wgt_9_160, // sfix19_En18 
  input [18:0] Wgt_9_161, // sfix19_En18 
  input [18:0] Wgt_9_162, // sfix19_En18 
  input [18:0] Wgt_9_163, // sfix19_En18 
  input [18:0] Wgt_9_164, // sfix19_En18 
  input [18:0] Wgt_9_165, // sfix19_En18 
  input [18:0] Wgt_9_166, // sfix19_En18 
  input [18:0] Wgt_9_167, // sfix19_En18 
  input [18:0] Wgt_9_168, // sfix19_En18 
  input [18:0] Wgt_9_169, // sfix19_En18 
  input [18:0] Wgt_9_170, // sfix19_En18 
  input [18:0] Wgt_9_171, // sfix19_En18 
  input [18:0] Wgt_9_172, // sfix19_En18 
  input [18:0] Wgt_9_173, // sfix19_En18 
  input [18:0] Wgt_9_174, // sfix19_En18 
  input [18:0] Wgt_9_175, // sfix19_En18 
  input [18:0] Wgt_9_176, // sfix19_En18 
  input [18:0] Wgt_9_177, // sfix19_En18 
  input [18:0] Wgt_9_178, // sfix19_En18 
  input [18:0] Wgt_9_179, // sfix19_En18 
  input [18:0] Wgt_9_180, // sfix19_En18 
  input [18:0] Wgt_9_181, // sfix19_En18 
  input [18:0] Wgt_9_182, // sfix19_En18 
  input [18:0] Wgt_9_183, // sfix19_En18 
  input [18:0] Wgt_9_184, // sfix19_En18 
  input [18:0] Wgt_9_185, // sfix19_En18 
  input [18:0] Wgt_9_186, // sfix19_En18 
  input [18:0] Wgt_9_187, // sfix19_En18 
  input [18:0] Wgt_9_188, // sfix19_En18 
  input [18:0] Wgt_9_189, // sfix19_En18 
  input [18:0] Wgt_9_190, // sfix19_En18 
  input [18:0] Wgt_9_191, // sfix19_En18 
  input [18:0] Wgt_9_192, // sfix19_En18 
  input [18:0] Wgt_9_193, // sfix19_En18 
  input [18:0] Wgt_9_194, // sfix19_En18 
  input [18:0] Wgt_9_195, // sfix19_En18 
  input [18:0] Wgt_9_196, // sfix19_En18 
  input [18:0] Wgt_9_197, // sfix19_En18 
  input [18:0] Wgt_9_198, // sfix19_En18 
  input [18:0] Wgt_9_199, // sfix19_En18 
  input [18:0] Wgt_9_200, // sfix19_En18 
  input [18:0] Wgt_9_201, // sfix19_En18 
  input [18:0] Wgt_9_202, // sfix19_En18 
  input [18:0] Wgt_9_203, // sfix19_En18 
  input [18:0] Wgt_9_204, // sfix19_En18 
  input [18:0] Wgt_9_205, // sfix19_En18 
  input [18:0] Wgt_9_206, // sfix19_En18 
  input [18:0] Wgt_9_207, // sfix19_En18 
  input [18:0] Wgt_9_208, // sfix19_En18 
  input [18:0] Wgt_9_209, // sfix19_En18 
  input [18:0] Wgt_9_210, // sfix19_En18 
  input [18:0] Wgt_9_211, // sfix19_En18 
  input [18:0] Wgt_9_212, // sfix19_En18 
  input [18:0] Wgt_9_213, // sfix19_En18 
  input [18:0] Wgt_9_214, // sfix19_En18 
  input [18:0] Wgt_9_215, // sfix19_En18 
  input [18:0] Wgt_9_216, // sfix19_En18 
  input [18:0] Wgt_9_217, // sfix19_En18 
  input [18:0] Wgt_9_218, // sfix19_En18 
  input [18:0] Wgt_9_219, // sfix19_En18 
  input [18:0] Wgt_9_220, // sfix19_En18 
  input [18:0] Wgt_9_221, // sfix19_En18 
  input [18:0] Wgt_9_222, // sfix19_En18 
  input [18:0] Wgt_9_223, // sfix19_En18 
  input [18:0] Wgt_9_224, // sfix19_En18 
  input [18:0] Wgt_9_225, // sfix19_En18 
  input [18:0] Wgt_9_226, // sfix19_En18 
  input [18:0] Wgt_9_227, // sfix19_En18 
  input [18:0] Wgt_9_228, // sfix19_En18 
  input [18:0] Wgt_9_229, // sfix19_En18 
  input [18:0] Wgt_9_230, // sfix19_En18 
  input [18:0] Wgt_9_231, // sfix19_En18 
  input [18:0] Wgt_9_232, // sfix19_En18 
  input [18:0] Wgt_9_233, // sfix19_En18 
  input [18:0] Wgt_9_234, // sfix19_En18 
  input [18:0] Wgt_9_235, // sfix19_En18 
  input [18:0] Wgt_9_236, // sfix19_En18 
  input [18:0] Wgt_9_237, // sfix19_En18 
  input [18:0] Wgt_9_238, // sfix19_En18 
  input [18:0] Wgt_9_239, // sfix19_En18 
  input [18:0] Wgt_9_240, // sfix19_En18 
  input [18:0] Wgt_9_241, // sfix19_En18 
  input [18:0] Wgt_9_242, // sfix19_En18 
  input [18:0] Wgt_9_243, // sfix19_En18 
  input [18:0] Wgt_9_244, // sfix19_En18 
  input [18:0] Wgt_9_245, // sfix19_En18 
  input [18:0] Wgt_9_246, // sfix19_En18 
  input [18:0] Wgt_9_247, // sfix19_En18 
  input [18:0] Wgt_9_248, // sfix19_En18 
  input [18:0] Wgt_9_249, // sfix19_En18 
  input [18:0] Wgt_9_250, // sfix19_En18 
  input [18:0] Wgt_9_251, // sfix19_En18 
  input [18:0] Wgt_9_252, // sfix19_En18 
  input [18:0] Wgt_9_253, // sfix19_En18 
  input [18:0] Wgt_9_254, // sfix19_En18 
  input [18:0] Wgt_9_255, // sfix19_En18 
  input [18:0] Wgt_9_256, // sfix19_En18 
  input [18:0] Wgt_9_257, // sfix19_En18 
  input [18:0] Wgt_9_258, // sfix19_En18 
  input [18:0] Wgt_9_259, // sfix19_En18 
  input [18:0] Wgt_9_260, // sfix19_En18 
  input [18:0] Wgt_9_261, // sfix19_En18 
  input [18:0] Wgt_9_262, // sfix19_En18 
  input [18:0] Wgt_9_263, // sfix19_En18 
  input [18:0] Wgt_9_264, // sfix19_En18 
  input [18:0] Wgt_9_265, // sfix19_En18 
  input [18:0] Wgt_9_266, // sfix19_En18 
  input [18:0] Wgt_9_267, // sfix19_En18 
  input [18:0] Wgt_9_268, // sfix19_En18 
  input [18:0] Wgt_9_269, // sfix19_En18 
  input [18:0] Wgt_9_270, // sfix19_En18 
  input [18:0] Wgt_9_271, // sfix19_En18 
  input [18:0] Wgt_9_272, // sfix19_En18 
  input [18:0] Wgt_9_273, // sfix19_En18 
  input [18:0] Wgt_9_274, // sfix19_En18 
  input [18:0] Wgt_9_275, // sfix19_En18 
  input [18:0] Wgt_9_276, // sfix19_En18 
  input [18:0] Wgt_9_277, // sfix19_En18 
  input [18:0] Wgt_9_278, // sfix19_En18 
  input [18:0] Wgt_9_279, // sfix19_En18 
  input [18:0] Wgt_9_280, // sfix19_En18 
  input [18:0] Wgt_9_281, // sfix19_En18 
  input [18:0] Wgt_9_282, // sfix19_En18 
  input [18:0] Wgt_9_283, // sfix19_En18 
  input [18:0] Wgt_9_284, // sfix19_En18 
  input [18:0] Wgt_9_285, // sfix19_En18 
  input [18:0] Wgt_9_286, // sfix19_En18 
  input [18:0] Wgt_9_287, // sfix19_En18 
  input [18:0] Wgt_9_288, // sfix19_En18 
  input [18:0] Wgt_9_289, // sfix19_En18 
  input [18:0] Wgt_9_290, // sfix19_En18 
  input [18:0] Wgt_9_291, // sfix19_En18 
  input [18:0] Wgt_9_292, // sfix19_En18 
  input [18:0] Wgt_9_293, // sfix19_En18 
  input [18:0] Wgt_9_294, // sfix19_En18 
  input [18:0] Wgt_9_295, // sfix19_En18 
  input [18:0] Wgt_9_296, // sfix19_En18 
  input [18:0] Wgt_9_297, // sfix19_En18 
  input [18:0] Wgt_9_298, // sfix19_En18 
  input [18:0] Wgt_9_299, // sfix19_En18 
  input [18:0] Wgt_9_300, // sfix19_En18 
  input [18:0] Wgt_9_301, // sfix19_En18 
  input [18:0] Wgt_9_302, // sfix19_En18 
  input [18:0] Wgt_9_303, // sfix19_En18 
  input [18:0] Wgt_9_304, // sfix19_En18 
  input [18:0] Wgt_9_305, // sfix19_En18 
  input [18:0] Wgt_9_306, // sfix19_En18 
  input [18:0] Wgt_9_307, // sfix19_En18 
  input [18:0] Wgt_9_308, // sfix19_En18 
  input [18:0] Wgt_9_309, // sfix19_En18 
  input [18:0] Wgt_9_310, // sfix19_En18 
  input [18:0] Wgt_9_311, // sfix19_En18 
  input [18:0] Wgt_9_312, // sfix19_En18 
  input [18:0] Wgt_9_313, // sfix19_En18 
  input [18:0] Wgt_9_314, // sfix19_En18 
  input [18:0] Wgt_9_315, // sfix19_En18 
  input [18:0] Wgt_9_316, // sfix19_En18 
  input [18:0] Wgt_9_317, // sfix19_En18 
  input [18:0] Wgt_9_318, // sfix19_En18 
  input [18:0] Wgt_9_319, // sfix19_En18 
  input [18:0] Wgt_9_320, // sfix19_En18 
  input [18:0] Wgt_9_321, // sfix19_En18 
  input [18:0] Wgt_9_322, // sfix19_En18 
  input [18:0] Wgt_9_323, // sfix19_En18 
  input [18:0] Wgt_9_324, // sfix19_En18 
  input [18:0] Wgt_9_325, // sfix19_En18 
  input [18:0] Wgt_9_326, // sfix19_En18 
  input [18:0] Wgt_9_327, // sfix19_En18 
  input [18:0] Wgt_9_328, // sfix19_En18 
  input [18:0] Wgt_9_329, // sfix19_En18 
  input [18:0] Wgt_9_330, // sfix19_En18 
  input [18:0] Wgt_9_331, // sfix19_En18 
  input [18:0] Wgt_9_332, // sfix19_En18 
  input [18:0] Wgt_9_333, // sfix19_En18 
  input [18:0] Wgt_9_334, // sfix19_En18 
  input [18:0] Wgt_9_335, // sfix19_En18 
  input [18:0] Wgt_9_336, // sfix19_En18 
  input [18:0] Wgt_9_337, // sfix19_En18 
  input [18:0] Wgt_9_338, // sfix19_En18 
  input [18:0] Wgt_9_339, // sfix19_En18 
  input [18:0] Wgt_9_340, // sfix19_En18 
  input [18:0] Wgt_9_341, // sfix19_En18 
  input [18:0] Wgt_9_342, // sfix19_En18 
  input [18:0] Wgt_9_343, // sfix19_En18 
  input [18:0] Wgt_9_344, // sfix19_En18 
  input [18:0] Wgt_9_345, // sfix19_En18 
  input [18:0] Wgt_9_346, // sfix19_En18 
  input [18:0] Wgt_9_347, // sfix19_En18 
  input [18:0] Wgt_9_348, // sfix19_En18 
  input [18:0] Wgt_9_349, // sfix19_En18 
  input [18:0] Wgt_9_350, // sfix19_En18 
  input [18:0] Wgt_9_351, // sfix19_En18 
  input [18:0] Wgt_9_352, // sfix19_En18 
  input [18:0] Wgt_9_353, // sfix19_En18 
  input [18:0] Wgt_9_354, // sfix19_En18 
  input [18:0] Wgt_9_355, // sfix19_En18 
  input [18:0] Wgt_9_356, // sfix19_En18 
  input [18:0] Wgt_9_357, // sfix19_En18 
  input [18:0] Wgt_9_358, // sfix19_En18 
  input [18:0] Wgt_9_359, // sfix19_En18 
  input [18:0] Wgt_9_360, // sfix19_En18 
  input [18:0] Wgt_9_361, // sfix19_En18 
  input [18:0] Wgt_9_362, // sfix19_En18 
  input [18:0] Wgt_9_363, // sfix19_En18 
  input [18:0] Wgt_9_364, // sfix19_En18 
  input [18:0] Wgt_9_365, // sfix19_En18 
  input [18:0] Wgt_9_366, // sfix19_En18 
  input [18:0] Wgt_9_367, // sfix19_En18 
  input [18:0] Wgt_9_368, // sfix19_En18 
  input [18:0] Wgt_9_369, // sfix19_En18 
  input [18:0] Wgt_9_370, // sfix19_En18 
  input [18:0] Wgt_9_371, // sfix19_En18 
  input [18:0] Wgt_9_372, // sfix19_En18 
  input [18:0] Wgt_9_373, // sfix19_En18 
  input [18:0] Wgt_9_374, // sfix19_En18 
  input [18:0] Wgt_9_375, // sfix19_En18 
  input [18:0] Wgt_9_376, // sfix19_En18 
  input [18:0] Wgt_9_377, // sfix19_En18 
  input [18:0] Wgt_9_378, // sfix19_En18 
  input [18:0] Wgt_9_379, // sfix19_En18 
  input [18:0] Wgt_9_380, // sfix19_En18 
  input [18:0] Wgt_9_381, // sfix19_En18 
  input [18:0] Wgt_9_382, // sfix19_En18 
  input [18:0] Wgt_9_383, // sfix19_En18 
  input [18:0] Wgt_9_384, // sfix19_En18 
  input [18:0] Wgt_9_385, // sfix19_En18 
  input [18:0] Wgt_9_386, // sfix19_En18 
  input [18:0] Wgt_9_387, // sfix19_En18 
  input [18:0] Wgt_9_388, // sfix19_En18 
  input [18:0] Wgt_9_389, // sfix19_En18 
  input [18:0] Wgt_9_390, // sfix19_En18 
  input [18:0] Wgt_9_391, // sfix19_En18 
  input [18:0] Wgt_9_392, // sfix19_En18 
  input [18:0] Wgt_9_393, // sfix19_En18 
  input [18:0] Wgt_9_394, // sfix19_En18 
  input [18:0] Wgt_9_395, // sfix19_En18 
  input [18:0] Wgt_9_396, // sfix19_En18 
  input [18:0] Wgt_9_397, // sfix19_En18 
  input [18:0] Wgt_9_398, // sfix19_En18 
  input [18:0] Wgt_9_399, // sfix19_En18 
  input [18:0] Wgt_9_400, // sfix19_En18 
  input [18:0] Wgt_9_401, // sfix19_En18 
  input [18:0] Wgt_9_402, // sfix19_En18 
  input [18:0] Wgt_9_403, // sfix19_En18 
  input [18:0] Wgt_9_404, // sfix19_En18 
  input [18:0] Wgt_9_405, // sfix19_En18 
  input [18:0] Wgt_9_406, // sfix19_En18 
  input [18:0] Wgt_9_407, // sfix19_En18 
  input [18:0] Wgt_9_408, // sfix19_En18 
  input [18:0] Wgt_9_409, // sfix19_En18 
  input [18:0] Wgt_9_410, // sfix19_En18 
  input [18:0] Wgt_9_411, // sfix19_En18 
  input [18:0] Wgt_9_412, // sfix19_En18 
  input [18:0] Wgt_9_413, // sfix19_En18 
  input [18:0] Wgt_9_414, // sfix19_En18 
  input [18:0] Wgt_9_415, // sfix19_En18 
  input [18:0] Wgt_9_416, // sfix19_En18 
  input [18:0] Wgt_9_417, // sfix19_En18 
  input [18:0] Wgt_9_418, // sfix19_En18 
  input [18:0] Wgt_9_419, // sfix19_En18 
  input [18:0] Wgt_9_420, // sfix19_En18 
  input [18:0] Wgt_9_421, // sfix19_En18 
  input [18:0] Wgt_9_422, // sfix19_En18 
  input [18:0] Wgt_9_423, // sfix19_En18 
  input [18:0] Wgt_9_424, // sfix19_En18 
  input [18:0] Wgt_9_425, // sfix19_En18 
  input [18:0] Wgt_9_426, // sfix19_En18 
  input [18:0] Wgt_9_427, // sfix19_En18 
  input [18:0] Wgt_9_428, // sfix19_En18 
  input [18:0] Wgt_9_429, // sfix19_En18 
  input [18:0] Wgt_9_430, // sfix19_En18 
  input [18:0] Wgt_9_431, // sfix19_En18 
  input [18:0] Wgt_9_432, // sfix19_En18 
  input [18:0] Wgt_9_433, // sfix19_En18 
  input [18:0] Wgt_9_434, // sfix19_En18 
  input [18:0] Wgt_9_435, // sfix19_En18 
  input [18:0] Wgt_9_436, // sfix19_En18 
  input [18:0] Wgt_9_437, // sfix19_En18 
  input [18:0] Wgt_9_438, // sfix19_En18 
  input [18:0] Wgt_9_439, // sfix19_En18 
  input [18:0] Wgt_9_440, // sfix19_En18 
  input [18:0] Wgt_9_441, // sfix19_En18 
  input [18:0] Wgt_9_442, // sfix19_En18 
  input [18:0] Wgt_9_443, // sfix19_En18 
  input [18:0] Wgt_9_444, // sfix19_En18 
  input [18:0] Wgt_9_445, // sfix19_En18 
  input [18:0] Wgt_9_446, // sfix19_En18 
  input [18:0] Wgt_9_447, // sfix19_En18 
  input [18:0] Wgt_9_448, // sfix19_En18 
  input [18:0] Wgt_9_449, // sfix19_En18 
  input [18:0] Wgt_9_450, // sfix19_En18 
  input [18:0] Wgt_9_451, // sfix19_En18 
  input [18:0] Wgt_9_452, // sfix19_En18 
  input [18:0] Wgt_9_453, // sfix19_En18 
  input [18:0] Wgt_9_454, // sfix19_En18 
  input [18:0] Wgt_9_455, // sfix19_En18 
  input [18:0] Wgt_9_456, // sfix19_En18 
  input [18:0] Wgt_9_457, // sfix19_En18 
  input [18:0] Wgt_9_458, // sfix19_En18 
  input [18:0] Wgt_9_459, // sfix19_En18 
  input [18:0] Wgt_9_460, // sfix19_En18 
  input [18:0] Wgt_9_461, // sfix19_En18 
  input [18:0] Wgt_9_462, // sfix19_En18 
  input [18:0] Wgt_9_463, // sfix19_En18 
  input [18:0] Wgt_9_464, // sfix19_En18 
  input [18:0] Wgt_9_465, // sfix19_En18 
  input [18:0] Wgt_9_466, // sfix19_En18 
  input [18:0] Wgt_9_467, // sfix19_En18 
  input [18:0] Wgt_9_468, // sfix19_En18 
  input [18:0] Wgt_9_469, // sfix19_En18 
  input [18:0] Wgt_9_470, // sfix19_En18 
  input [18:0] Wgt_9_471, // sfix19_En18 
  input [18:0] Wgt_9_472, // sfix19_En18 
  input [18:0] Wgt_9_473, // sfix19_En18 
  input [18:0] Wgt_9_474, // sfix19_En18 
  input [18:0] Wgt_9_475, // sfix19_En18 
  input [18:0] Wgt_9_476, // sfix19_En18 
  input [18:0] Wgt_9_477, // sfix19_En18 
  input [18:0] Wgt_9_478, // sfix19_En18 
  input [18:0] Wgt_9_479, // sfix19_En18 
  input [18:0] Wgt_9_480, // sfix19_En18 
  input [18:0] Wgt_9_481, // sfix19_En18 
  input [18:0] Wgt_9_482, // sfix19_En18 
  input [18:0] Wgt_9_483, // sfix19_En18 
  input [18:0] Wgt_9_484, // sfix19_En18 
  input [18:0] Wgt_9_485, // sfix19_En18 
  input [18:0] Wgt_9_486, // sfix19_En18 
  input [18:0] Wgt_9_487, // sfix19_En18 
  input [18:0] Wgt_9_488, // sfix19_En18 
  input [18:0] Wgt_9_489, // sfix19_En18 
  input [18:0] Wgt_9_490, // sfix19_En18 
  input [18:0] Wgt_9_491, // sfix19_En18 
  input [18:0] Wgt_9_492, // sfix19_En18 
  input [18:0] Wgt_9_493, // sfix19_En18 
  input [18:0] Wgt_9_494, // sfix19_En18 
  input [18:0] Wgt_9_495, // sfix19_En18 
  input [18:0] Wgt_9_496, // sfix19_En18 
  input [18:0] Wgt_9_497, // sfix19_En18 
  input [18:0] Wgt_9_498, // sfix19_En18 
  input [18:0] Wgt_9_499, // sfix19_En18 
  input [18:0] Wgt_9_500, // sfix19_En18 
  input [18:0] Wgt_9_501, // sfix19_En18 
  input [18:0] Wgt_9_502, // sfix19_En18 
  input [18:0] Wgt_9_503, // sfix19_En18 
  input [18:0] Wgt_9_504, // sfix19_En18 
  input [18:0] Wgt_9_505, // sfix19_En18 
  input [18:0] Wgt_9_506, // sfix19_En18 
  input [18:0] Wgt_9_507, // sfix19_En18 
  input [18:0] Wgt_9_508, // sfix19_En18 
  input [18:0] Wgt_9_509, // sfix19_En18 
  input [18:0] Wgt_9_510, // sfix19_En18 
  input [18:0] Wgt_9_511, // sfix19_En18 
  input [18:0] Wgt_9_512, // sfix19_En18 
  input [18:0] Wgt_9_513, // sfix19_En18 
  input [18:0] Wgt_9_514, // sfix19_En18 
  input [18:0] Wgt_9_515, // sfix19_En18 
  input [18:0] Wgt_9_516, // sfix19_En18 
  input [18:0] Wgt_9_517, // sfix19_En18 
  input [18:0] Wgt_9_518, // sfix19_En18 
  input [18:0] Wgt_9_519, // sfix19_En18 
  input [18:0] Wgt_9_520, // sfix19_En18 
  input [18:0] Wgt_9_521, // sfix19_En18 
  input [18:0] Wgt_9_522, // sfix19_En18 
  input [18:0] Wgt_9_523, // sfix19_En18 
  input [18:0] Wgt_9_524, // sfix19_En18 
  input [18:0] Wgt_9_525, // sfix19_En18 
  input [18:0] Wgt_9_526, // sfix19_En18 
  input [18:0] Wgt_9_527, // sfix19_En18 
  input [18:0] Wgt_9_528, // sfix19_En18 
  input [18:0] Wgt_9_529, // sfix19_En18 
  input [18:0] Wgt_9_530, // sfix19_En18 
  input [18:0] Wgt_9_531, // sfix19_En18 
  input [18:0] Wgt_9_532, // sfix19_En18 
  input [18:0] Wgt_9_533, // sfix19_En18 
  input [18:0] Wgt_9_534, // sfix19_En18 
  input [18:0] Wgt_9_535, // sfix19_En18 
  input [18:0] Wgt_9_536, // sfix19_En18 
  input [18:0] Wgt_9_537, // sfix19_En18 
  input [18:0] Wgt_9_538, // sfix19_En18 
  input [18:0] Wgt_9_539, // sfix19_En18 
  input [18:0] Wgt_9_540, // sfix19_En18 
  input [18:0] Wgt_9_541, // sfix19_En18 
  input [18:0] Wgt_9_542, // sfix19_En18 
  input [18:0] Wgt_9_543, // sfix19_En18 
  input [18:0] Wgt_9_544, // sfix19_En18 
  input [18:0] Wgt_9_545, // sfix19_En18 
  input [18:0] Wgt_9_546, // sfix19_En18 
  input [18:0] Wgt_9_547, // sfix19_En18 
  input [18:0] Wgt_9_548, // sfix19_En18 
  input [18:0] Wgt_9_549, // sfix19_En18 
  input [18:0] Wgt_9_550, // sfix19_En18 
  input [18:0] Wgt_9_551, // sfix19_En18 
  input [18:0] Wgt_9_552, // sfix19_En18 
  input [18:0] Wgt_9_553, // sfix19_En18 
  input [18:0] Wgt_9_554, // sfix19_En18 
  input [18:0] Wgt_9_555, // sfix19_En18 
  input [18:0] Wgt_9_556, // sfix19_En18 
  input [18:0] Wgt_9_557, // sfix19_En18 
  input [18:0] Wgt_9_558, // sfix19_En18 
  input [18:0] Wgt_9_559, // sfix19_En18 
  input [18:0] Wgt_9_560, // sfix19_En18 
  input [18:0] Wgt_9_561, // sfix19_En18 
  input [18:0] Wgt_9_562, // sfix19_En18 
  input [18:0] Wgt_9_563, // sfix19_En18 
  input [18:0] Wgt_9_564, // sfix19_En18 
  input [18:0] Wgt_9_565, // sfix19_En18 
  input [18:0] Wgt_9_566, // sfix19_En18 
  input [18:0] Wgt_9_567, // sfix19_En18 
  input [18:0] Wgt_9_568, // sfix19_En18 
  input [18:0] Wgt_9_569, // sfix19_En18 
  input [18:0] Wgt_9_570, // sfix19_En18 
  input [18:0] Wgt_9_571, // sfix19_En18 
  input [18:0] Wgt_9_572, // sfix19_En18 
  input [18:0] Wgt_9_573, // sfix19_En18 
  input [18:0] Wgt_9_574, // sfix19_En18 
  input [18:0] Wgt_9_575, // sfix19_En18 
  input [18:0] Wgt_9_576, // sfix19_En18 
  input [18:0] Wgt_9_577, // sfix19_En18 
  input [18:0] Wgt_9_578, // sfix19_En18 
  input [18:0] Wgt_9_579, // sfix19_En18 
  input [18:0] Wgt_9_580, // sfix19_En18 
  input [18:0] Wgt_9_581, // sfix19_En18 
  input [18:0] Wgt_9_582, // sfix19_En18 
  input [18:0] Wgt_9_583, // sfix19_En18 
  input [18:0] Wgt_9_584, // sfix19_En18 
  input [18:0] Wgt_9_585, // sfix19_En18 
  input [18:0] Wgt_9_586, // sfix19_En18 
  input [18:0] Wgt_9_587, // sfix19_En18 
  input [18:0] Wgt_9_588, // sfix19_En18 
  input [18:0] Wgt_9_589, // sfix19_En18 
  input [18:0] Wgt_9_590, // sfix19_En18 
  input [18:0] Wgt_9_591, // sfix19_En18 
  input [18:0] Wgt_9_592, // sfix19_En18 
  input [18:0] Wgt_9_593, // sfix19_En18 
  input [18:0] Wgt_9_594, // sfix19_En18 
  input [18:0] Wgt_9_595, // sfix19_En18 
  input [18:0] Wgt_9_596, // sfix19_En18 
  input [18:0] Wgt_9_597, // sfix19_En18 
  input [18:0] Wgt_9_598, // sfix19_En18 
  input [18:0] Wgt_9_599, // sfix19_En18 
  input [18:0] Wgt_9_600, // sfix19_En18 
  input [18:0] Wgt_9_601, // sfix19_En18 
  input [18:0] Wgt_9_602, // sfix19_En18 
  input [18:0] Wgt_9_603, // sfix19_En18 
  input [18:0] Wgt_9_604, // sfix19_En18 
  input [18:0] Wgt_9_605, // sfix19_En18 
  input [18:0] Wgt_9_606, // sfix19_En18 
  input [18:0] Wgt_9_607, // sfix19_En18 
  input [18:0] Wgt_9_608, // sfix19_En18 
  input [18:0] Wgt_9_609, // sfix19_En18 
  input [18:0] Wgt_9_610, // sfix19_En18 
  input [18:0] Wgt_9_611, // sfix19_En18 
  input [18:0] Wgt_9_612, // sfix19_En18 
  input [18:0] Wgt_9_613, // sfix19_En18 
  input [18:0] Wgt_9_614, // sfix19_En18 
  input [18:0] Wgt_9_615, // sfix19_En18 
  input [18:0] Wgt_9_616, // sfix19_En18 
  input [18:0] Wgt_9_617, // sfix19_En18 
  input [18:0] Wgt_9_618, // sfix19_En18 
  input [18:0] Wgt_9_619, // sfix19_En18 
  input [18:0] Wgt_9_620, // sfix19_En18 
  input [18:0] Wgt_9_621, // sfix19_En18 
  input [18:0] Wgt_9_622, // sfix19_En18 
  input [18:0] Wgt_9_623, // sfix19_En18 
  input [18:0] Wgt_9_624, // sfix19_En18 
  input [18:0] Wgt_9_625, // sfix19_En18 
  input [18:0] Wgt_9_626, // sfix19_En18 
  input [18:0] Wgt_9_627, // sfix19_En18 
  input [18:0] Wgt_9_628, // sfix19_En18 
  input [18:0] Wgt_9_629, // sfix19_En18 
  input [18:0] Wgt_9_630, // sfix19_En18 
  input [18:0] Wgt_9_631, // sfix19_En18 
  input [18:0] Wgt_9_632, // sfix19_En18 
  input [18:0] Wgt_9_633, // sfix19_En18 
  input [18:0] Wgt_9_634, // sfix19_En18 
  input [18:0] Wgt_9_635, // sfix19_En18 
  input [18:0] Wgt_9_636, // sfix19_En18 
  input [18:0] Wgt_9_637, // sfix19_En18 
  input [18:0] Wgt_9_638, // sfix19_En18 
  input [18:0] Wgt_9_639, // sfix19_En18 
  input [18:0] Wgt_9_640, // sfix19_En18 
  input [18:0] Wgt_9_641, // sfix19_En18 
  input [18:0] Wgt_9_642, // sfix19_En18 
  input [18:0] Wgt_9_643, // sfix19_En18 
  input [18:0] Wgt_9_644, // sfix19_En18 
  input [18:0] Wgt_9_645, // sfix19_En18 
  input [18:0] Wgt_9_646, // sfix19_En18 
  input [18:0] Wgt_9_647, // sfix19_En18 
  input [18:0] Wgt_9_648, // sfix19_En18 
  input [18:0] Wgt_9_649, // sfix19_En18 
  input [18:0] Wgt_9_650, // sfix19_En18 
  input [18:0] Wgt_9_651, // sfix19_En18 
  input [18:0] Wgt_9_652, // sfix19_En18 
  input [18:0] Wgt_9_653, // sfix19_En18 
  input [18:0] Wgt_9_654, // sfix19_En18 
  input [18:0] Wgt_9_655, // sfix19_En18 
  input [18:0] Wgt_9_656, // sfix19_En18 
  input [18:0] Wgt_9_657, // sfix19_En18 
  input [18:0] Wgt_9_658, // sfix19_En18 
  input [18:0] Wgt_9_659, // sfix19_En18 
  input [18:0] Wgt_9_660, // sfix19_En18 
  input [18:0] Wgt_9_661, // sfix19_En18 
  input [18:0] Wgt_9_662, // sfix19_En18 
  input [18:0] Wgt_9_663, // sfix19_En18 
  input [18:0] Wgt_9_664, // sfix19_En18 
  input [18:0] Wgt_9_665, // sfix19_En18 
  input [18:0] Wgt_9_666, // sfix19_En18 
  input [18:0] Wgt_9_667, // sfix19_En18 
  input [18:0] Wgt_9_668, // sfix19_En18 
  input [18:0] Wgt_9_669, // sfix19_En18 
  input [18:0] Wgt_9_670, // sfix19_En18 
  input [18:0] Wgt_9_671, // sfix19_En18 
  input [18:0] Wgt_9_672, // sfix19_En18 
  input [18:0] Wgt_9_673, // sfix19_En18 
  input [18:0] Wgt_9_674, // sfix19_En18 
  input [18:0] Wgt_9_675, // sfix19_En18 
  input [18:0] Wgt_9_676, // sfix19_En18 
  input [18:0] Wgt_9_677, // sfix19_En18 
  input [18:0] Wgt_9_678, // sfix19_En18 
  input [18:0] Wgt_9_679, // sfix19_En18 
  input [18:0] Wgt_9_680, // sfix19_En18 
  input [18:0] Wgt_9_681, // sfix19_En18 
  input [18:0] Wgt_9_682, // sfix19_En18 
  input [18:0] Wgt_9_683, // sfix19_En18 
  input [18:0] Wgt_9_684, // sfix19_En18 
  input [18:0] Wgt_9_685, // sfix19_En18 
  input [18:0] Wgt_9_686, // sfix19_En18 
  input [18:0] Wgt_9_687, // sfix19_En18 
  input [18:0] Wgt_9_688, // sfix19_En18 
  input [18:0] Wgt_9_689, // sfix19_En18 
  input [18:0] Wgt_9_690, // sfix19_En18 
  input [18:0] Wgt_9_691, // sfix19_En18 
  input [18:0] Wgt_9_692, // sfix19_En18 
  input [18:0] Wgt_9_693, // sfix19_En18 
  input [18:0] Wgt_9_694, // sfix19_En18 
  input [18:0] Wgt_9_695, // sfix19_En18 
  input [18:0] Wgt_9_696, // sfix19_En18 
  input [18:0] Wgt_9_697, // sfix19_En18 
  input [18:0] Wgt_9_698, // sfix19_En18 
  input [18:0] Wgt_9_699, // sfix19_En18 
  input [18:0] Wgt_9_700, // sfix19_En18 
  input [18:0] Wgt_9_701, // sfix19_En18 
  input [18:0] Wgt_9_702, // sfix19_En18 
  input [18:0] Wgt_9_703, // sfix19_En18 
  input [18:0] Wgt_9_704, // sfix19_En18 
  input [18:0] Wgt_9_705, // sfix19_En18 
  input [18:0] Wgt_9_706, // sfix19_En18 
  input [18:0] Wgt_9_707, // sfix19_En18 
  input [18:0] Wgt_9_708, // sfix19_En18 
  input [18:0] Wgt_9_709, // sfix19_En18 
  input [18:0] Wgt_9_710, // sfix19_En18 
  input [18:0] Wgt_9_711, // sfix19_En18 
  input [18:0] Wgt_9_712, // sfix19_En18 
  input [18:0] Wgt_9_713, // sfix19_En18 
  input [18:0] Wgt_9_714, // sfix19_En18 
  input [18:0] Wgt_9_715, // sfix19_En18 
  input [18:0] Wgt_9_716, // sfix19_En18 
  input [18:0] Wgt_9_717, // sfix19_En18 
  input [18:0] Wgt_9_718, // sfix19_En18 
  input [18:0] Wgt_9_719, // sfix19_En18 
  input [18:0] Wgt_9_720, // sfix19_En18 
  input [18:0] Wgt_9_721, // sfix19_En18 
  input [18:0] Wgt_9_722, // sfix19_En18 
  input [18:0] Wgt_9_723, // sfix19_En18 
  input [18:0] Wgt_9_724, // sfix19_En18 
  input [18:0] Wgt_9_725, // sfix19_En18 
  input [18:0] Wgt_9_726, // sfix19_En18 
  input [18:0] Wgt_9_727, // sfix19_En18 
  input [18:0] Wgt_9_728, // sfix19_En18 
  input [18:0] Wgt_9_729, // sfix19_En18 
  input [18:0] Wgt_9_730, // sfix19_En18 
  input [18:0] Wgt_9_731, // sfix19_En18 
  input [18:0] Wgt_9_732, // sfix19_En18 
  input [18:0] Wgt_9_733, // sfix19_En18 
  input [18:0] Wgt_9_734, // sfix19_En18 
  input [18:0] Wgt_9_735, // sfix19_En18 
  input [18:0] Wgt_9_736, // sfix19_En18 
  input [18:0] Wgt_9_737, // sfix19_En18 
  input [18:0] Wgt_9_738, // sfix19_En18 
  input [18:0] Wgt_9_739, // sfix19_En18 
  input [18:0] Wgt_9_740, // sfix19_En18 
  input [18:0] Wgt_9_741, // sfix19_En18 
  input [18:0] Wgt_9_742, // sfix19_En18 
  input [18:0] Wgt_9_743, // sfix19_En18 
  input [18:0] Wgt_9_744, // sfix19_En18 
  input [18:0] Wgt_9_745, // sfix19_En18 
  input [18:0] Wgt_9_746, // sfix19_En18 
  input [18:0] Wgt_9_747, // sfix19_En18 
  input [18:0] Wgt_9_748, // sfix19_En18 
  input [18:0] Wgt_9_749, // sfix19_En18 
  input [18:0] Wgt_9_750, // sfix19_En18 
  input [18:0] Wgt_9_751, // sfix19_En18 
  input [18:0] Wgt_9_752, // sfix19_En18 
  input [18:0] Wgt_9_753, // sfix19_En18 
  input [18:0] Wgt_9_754, // sfix19_En18 
  input [18:0] Wgt_9_755, // sfix19_En18 
  input [18:0] Wgt_9_756, // sfix19_En18 
  input [18:0] Wgt_9_757, // sfix19_En18 
  input [18:0] Wgt_9_758, // sfix19_En18 
  input [18:0] Wgt_9_759, // sfix19_En18 
  input [18:0] Wgt_9_760, // sfix19_En18 
  input [18:0] Wgt_9_761, // sfix19_En18 
  input [18:0] Wgt_9_762, // sfix19_En18 
  input [18:0] Wgt_9_763, // sfix19_En18 
  input [18:0] Wgt_9_764, // sfix19_En18 
  input [18:0] Wgt_9_765, // sfix19_En18 
  input [18:0] Wgt_9_766, // sfix19_En18 
  input [18:0] Wgt_9_767, // sfix19_En18 
  input [18:0] Wgt_9_768, // sfix19_En18 
  input [18:0] Wgt_9_769, // sfix19_En18 
  input [18:0] Wgt_9_770, // sfix19_En18 
  input [18:0] Wgt_9_771, // sfix19_En18 
  input [18:0] Wgt_9_772, // sfix19_En18 
  input [18:0] Wgt_9_773, // sfix19_En18 
  input [18:0] Wgt_9_774, // sfix19_En18 
  input [18:0] Wgt_9_775, // sfix19_En18 
  input [18:0] Wgt_9_776, // sfix19_En18 
  input [18:0] Wgt_9_777, // sfix19_En18 
  input [18:0] Wgt_9_778, // sfix19_En18 
  input [18:0] Wgt_9_779, // sfix19_En18 
  input [18:0] Wgt_9_780, // sfix19_En18 
  input [18:0] Wgt_9_781, // sfix19_En18 
  input [18:0] Wgt_9_782, // sfix19_En18 
  input [18:0] Wgt_9_783, // sfix19_En18 
  input [18:0] Wgt_9_784, // sfix19_En18 
  input [9:0] Pix_0, // sfix10_En0 
 input [9:0] Pix_1, // sfix10_En0 
 input [9:0] Pix_2, // sfix10_En0 
 input [9:0] Pix_3, // sfix10_En0 
 input [9:0] Pix_4, // sfix10_En0 
 input [9:0] Pix_5, // sfix10_En0 
 input [9:0] Pix_6, // sfix10_En0 
 input [9:0] Pix_7, // sfix10_En0 
 input [9:0] Pix_8, // sfix10_En0 
 input [9:0] Pix_9, // sfix10_En0 
 input [9:0] Pix_10, // sfix10_En0 
 input [9:0] Pix_11, // sfix10_En0 
 input [9:0] Pix_12, // sfix10_En0 
 input [9:0] Pix_13, // sfix10_En0 
 input [9:0] Pix_14, // sfix10_En0 
 input [9:0] Pix_15, // sfix10_En0 
 input [9:0] Pix_16, // sfix10_En0 
 input [9:0] Pix_17, // sfix10_En0 
 input [9:0] Pix_18, // sfix10_En0 
 input [9:0] Pix_19, // sfix10_En0 
 input [9:0] Pix_20, // sfix10_En0 
 input [9:0] Pix_21, // sfix10_En0 
 input [9:0] Pix_22, // sfix10_En0 
 input [9:0] Pix_23, // sfix10_En0 
 input [9:0] Pix_24, // sfix10_En0 
 input [9:0] Pix_25, // sfix10_En0 
 input [9:0] Pix_26, // sfix10_En0 
 input [9:0] Pix_27, // sfix10_En0 
 input [9:0] Pix_28, // sfix10_En0 
 input [9:0] Pix_29, // sfix10_En0 
 input [9:0] Pix_30, // sfix10_En0 
 input [9:0] Pix_31, // sfix10_En0 
 input [9:0] Pix_32, // sfix10_En0 
 input [9:0] Pix_33, // sfix10_En0 
 input [9:0] Pix_34, // sfix10_En0 
 input [9:0] Pix_35, // sfix10_En0 
 input [9:0] Pix_36, // sfix10_En0 
 input [9:0] Pix_37, // sfix10_En0 
 input [9:0] Pix_38, // sfix10_En0 
 input [9:0] Pix_39, // sfix10_En0 
 input [9:0] Pix_40, // sfix10_En0 
 input [9:0] Pix_41, // sfix10_En0 
 input [9:0] Pix_42, // sfix10_En0 
 input [9:0] Pix_43, // sfix10_En0 
 input [9:0] Pix_44, // sfix10_En0 
 input [9:0] Pix_45, // sfix10_En0 
 input [9:0] Pix_46, // sfix10_En0 
 input [9:0] Pix_47, // sfix10_En0 
 input [9:0] Pix_48, // sfix10_En0 
 input [9:0] Pix_49, // sfix10_En0 
 input [9:0] Pix_50, // sfix10_En0 
 input [9:0] Pix_51, // sfix10_En0 
 input [9:0] Pix_52, // sfix10_En0 
 input [9:0] Pix_53, // sfix10_En0 
 input [9:0] Pix_54, // sfix10_En0 
 input [9:0] Pix_55, // sfix10_En0 
 input [9:0] Pix_56, // sfix10_En0 
 input [9:0] Pix_57, // sfix10_En0 
 input [9:0] Pix_58, // sfix10_En0 
 input [9:0] Pix_59, // sfix10_En0 
 input [9:0] Pix_60, // sfix10_En0 
 input [9:0] Pix_61, // sfix10_En0 
 input [9:0] Pix_62, // sfix10_En0 
 input [9:0] Pix_63, // sfix10_En0 
 input [9:0] Pix_64, // sfix10_En0 
 input [9:0] Pix_65, // sfix10_En0 
 input [9:0] Pix_66, // sfix10_En0 
 input [9:0] Pix_67, // sfix10_En0 
 input [9:0] Pix_68, // sfix10_En0 
 input [9:0] Pix_69, // sfix10_En0 
 input [9:0] Pix_70, // sfix10_En0 
 input [9:0] Pix_71, // sfix10_En0 
 input [9:0] Pix_72, // sfix10_En0 
 input [9:0] Pix_73, // sfix10_En0 
 input [9:0] Pix_74, // sfix10_En0 
 input [9:0] Pix_75, // sfix10_En0 
 input [9:0] Pix_76, // sfix10_En0 
 input [9:0] Pix_77, // sfix10_En0 
 input [9:0] Pix_78, // sfix10_En0 
 input [9:0] Pix_79, // sfix10_En0 
 input [9:0] Pix_80, // sfix10_En0 
 input [9:0] Pix_81, // sfix10_En0 
 input [9:0] Pix_82, // sfix10_En0 
 input [9:0] Pix_83, // sfix10_En0 
 input [9:0] Pix_84, // sfix10_En0 
 input [9:0] Pix_85, // sfix10_En0 
 input [9:0] Pix_86, // sfix10_En0 
 input [9:0] Pix_87, // sfix10_En0 
 input [9:0] Pix_88, // sfix10_En0 
 input [9:0] Pix_89, // sfix10_En0 
 input [9:0] Pix_90, // sfix10_En0 
 input [9:0] Pix_91, // sfix10_En0 
 input [9:0] Pix_92, // sfix10_En0 
 input [9:0] Pix_93, // sfix10_En0 
 input [9:0] Pix_94, // sfix10_En0 
 input [9:0] Pix_95, // sfix10_En0 
 input [9:0] Pix_96, // sfix10_En0 
 input [9:0] Pix_97, // sfix10_En0 
 input [9:0] Pix_98, // sfix10_En0 
 input [9:0] Pix_99, // sfix10_En0 
 input [9:0] Pix_100, // sfix10_En0 
 input [9:0] Pix_101, // sfix10_En0 
 input [9:0] Pix_102, // sfix10_En0 
 input [9:0] Pix_103, // sfix10_En0 
 input [9:0] Pix_104, // sfix10_En0 
 input [9:0] Pix_105, // sfix10_En0 
 input [9:0] Pix_106, // sfix10_En0 
 input [9:0] Pix_107, // sfix10_En0 
 input [9:0] Pix_108, // sfix10_En0 
 input [9:0] Pix_109, // sfix10_En0 
 input [9:0] Pix_110, // sfix10_En0 
 input [9:0] Pix_111, // sfix10_En0 
 input [9:0] Pix_112, // sfix10_En0 
 input [9:0] Pix_113, // sfix10_En0 
 input [9:0] Pix_114, // sfix10_En0 
 input [9:0] Pix_115, // sfix10_En0 
 input [9:0] Pix_116, // sfix10_En0 
 input [9:0] Pix_117, // sfix10_En0 
 input [9:0] Pix_118, // sfix10_En0 
 input [9:0] Pix_119, // sfix10_En0 
 input [9:0] Pix_120, // sfix10_En0 
 input [9:0] Pix_121, // sfix10_En0 
 input [9:0] Pix_122, // sfix10_En0 
 input [9:0] Pix_123, // sfix10_En0 
 input [9:0] Pix_124, // sfix10_En0 
 input [9:0] Pix_125, // sfix10_En0 
 input [9:0] Pix_126, // sfix10_En0 
 input [9:0] Pix_127, // sfix10_En0 
 input [9:0] Pix_128, // sfix10_En0 
 input [9:0] Pix_129, // sfix10_En0 
 input [9:0] Pix_130, // sfix10_En0 
 input [9:0] Pix_131, // sfix10_En0 
 input [9:0] Pix_132, // sfix10_En0 
 input [9:0] Pix_133, // sfix10_En0 
 input [9:0] Pix_134, // sfix10_En0 
 input [9:0] Pix_135, // sfix10_En0 
 input [9:0] Pix_136, // sfix10_En0 
 input [9:0] Pix_137, // sfix10_En0 
 input [9:0] Pix_138, // sfix10_En0 
 input [9:0] Pix_139, // sfix10_En0 
 input [9:0] Pix_140, // sfix10_En0 
 input [9:0] Pix_141, // sfix10_En0 
 input [9:0] Pix_142, // sfix10_En0 
 input [9:0] Pix_143, // sfix10_En0 
 input [9:0] Pix_144, // sfix10_En0 
 input [9:0] Pix_145, // sfix10_En0 
 input [9:0] Pix_146, // sfix10_En0 
 input [9:0] Pix_147, // sfix10_En0 
 input [9:0] Pix_148, // sfix10_En0 
 input [9:0] Pix_149, // sfix10_En0 
 input [9:0] Pix_150, // sfix10_En0 
 input [9:0] Pix_151, // sfix10_En0 
 input [9:0] Pix_152, // sfix10_En0 
 input [9:0] Pix_153, // sfix10_En0 
 input [9:0] Pix_154, // sfix10_En0 
 input [9:0] Pix_155, // sfix10_En0 
 input [9:0] Pix_156, // sfix10_En0 
 input [9:0] Pix_157, // sfix10_En0 
 input [9:0] Pix_158, // sfix10_En0 
 input [9:0] Pix_159, // sfix10_En0 
 input [9:0] Pix_160, // sfix10_En0 
 input [9:0] Pix_161, // sfix10_En0 
 input [9:0] Pix_162, // sfix10_En0 
 input [9:0] Pix_163, // sfix10_En0 
 input [9:0] Pix_164, // sfix10_En0 
 input [9:0] Pix_165, // sfix10_En0 
 input [9:0] Pix_166, // sfix10_En0 
 input [9:0] Pix_167, // sfix10_En0 
 input [9:0] Pix_168, // sfix10_En0 
 input [9:0] Pix_169, // sfix10_En0 
 input [9:0] Pix_170, // sfix10_En0 
 input [9:0] Pix_171, // sfix10_En0 
 input [9:0] Pix_172, // sfix10_En0 
 input [9:0] Pix_173, // sfix10_En0 
 input [9:0] Pix_174, // sfix10_En0 
 input [9:0] Pix_175, // sfix10_En0 
 input [9:0] Pix_176, // sfix10_En0 
 input [9:0] Pix_177, // sfix10_En0 
 input [9:0] Pix_178, // sfix10_En0 
 input [9:0] Pix_179, // sfix10_En0 
 input [9:0] Pix_180, // sfix10_En0 
 input [9:0] Pix_181, // sfix10_En0 
 input [9:0] Pix_182, // sfix10_En0 
 input [9:0] Pix_183, // sfix10_En0 
 input [9:0] Pix_184, // sfix10_En0 
 input [9:0] Pix_185, // sfix10_En0 
 input [9:0] Pix_186, // sfix10_En0 
 input [9:0] Pix_187, // sfix10_En0 
 input [9:0] Pix_188, // sfix10_En0 
 input [9:0] Pix_189, // sfix10_En0 
 input [9:0] Pix_190, // sfix10_En0 
 input [9:0] Pix_191, // sfix10_En0 
 input [9:0] Pix_192, // sfix10_En0 
 input [9:0] Pix_193, // sfix10_En0 
 input [9:0] Pix_194, // sfix10_En0 
 input [9:0] Pix_195, // sfix10_En0 
 input [9:0] Pix_196, // sfix10_En0 
 input [9:0] Pix_197, // sfix10_En0 
 input [9:0] Pix_198, // sfix10_En0 
 input [9:0] Pix_199, // sfix10_En0 
 input [9:0] Pix_200, // sfix10_En0 
 input [9:0] Pix_201, // sfix10_En0 
 input [9:0] Pix_202, // sfix10_En0 
 input [9:0] Pix_203, // sfix10_En0 
 input [9:0] Pix_204, // sfix10_En0 
 input [9:0] Pix_205, // sfix10_En0 
 input [9:0] Pix_206, // sfix10_En0 
 input [9:0] Pix_207, // sfix10_En0 
 input [9:0] Pix_208, // sfix10_En0 
 input [9:0] Pix_209, // sfix10_En0 
 input [9:0] Pix_210, // sfix10_En0 
 input [9:0] Pix_211, // sfix10_En0 
 input [9:0] Pix_212, // sfix10_En0 
 input [9:0] Pix_213, // sfix10_En0 
 input [9:0] Pix_214, // sfix10_En0 
 input [9:0] Pix_215, // sfix10_En0 
 input [9:0] Pix_216, // sfix10_En0 
 input [9:0] Pix_217, // sfix10_En0 
 input [9:0] Pix_218, // sfix10_En0 
 input [9:0] Pix_219, // sfix10_En0 
 input [9:0] Pix_220, // sfix10_En0 
 input [9:0] Pix_221, // sfix10_En0 
 input [9:0] Pix_222, // sfix10_En0 
 input [9:0] Pix_223, // sfix10_En0 
 input [9:0] Pix_224, // sfix10_En0 
 input [9:0] Pix_225, // sfix10_En0 
 input [9:0] Pix_226, // sfix10_En0 
 input [9:0] Pix_227, // sfix10_En0 
 input [9:0] Pix_228, // sfix10_En0 
 input [9:0] Pix_229, // sfix10_En0 
 input [9:0] Pix_230, // sfix10_En0 
 input [9:0] Pix_231, // sfix10_En0 
 input [9:0] Pix_232, // sfix10_En0 
 input [9:0] Pix_233, // sfix10_En0 
 input [9:0] Pix_234, // sfix10_En0 
 input [9:0] Pix_235, // sfix10_En0 
 input [9:0] Pix_236, // sfix10_En0 
 input [9:0] Pix_237, // sfix10_En0 
 input [9:0] Pix_238, // sfix10_En0 
 input [9:0] Pix_239, // sfix10_En0 
 input [9:0] Pix_240, // sfix10_En0 
 input [9:0] Pix_241, // sfix10_En0 
 input [9:0] Pix_242, // sfix10_En0 
 input [9:0] Pix_243, // sfix10_En0 
 input [9:0] Pix_244, // sfix10_En0 
 input [9:0] Pix_245, // sfix10_En0 
 input [9:0] Pix_246, // sfix10_En0 
 input [9:0] Pix_247, // sfix10_En0 
 input [9:0] Pix_248, // sfix10_En0 
 input [9:0] Pix_249, // sfix10_En0 
 input [9:0] Pix_250, // sfix10_En0 
 input [9:0] Pix_251, // sfix10_En0 
 input [9:0] Pix_252, // sfix10_En0 
 input [9:0] Pix_253, // sfix10_En0 
 input [9:0] Pix_254, // sfix10_En0 
 input [9:0] Pix_255, // sfix10_En0 
 input [9:0] Pix_256, // sfix10_En0 
 input [9:0] Pix_257, // sfix10_En0 
 input [9:0] Pix_258, // sfix10_En0 
 input [9:0] Pix_259, // sfix10_En0 
 input [9:0] Pix_260, // sfix10_En0 
 input [9:0] Pix_261, // sfix10_En0 
 input [9:0] Pix_262, // sfix10_En0 
 input [9:0] Pix_263, // sfix10_En0 
 input [9:0] Pix_264, // sfix10_En0 
 input [9:0] Pix_265, // sfix10_En0 
 input [9:0] Pix_266, // sfix10_En0 
 input [9:0] Pix_267, // sfix10_En0 
 input [9:0] Pix_268, // sfix10_En0 
 input [9:0] Pix_269, // sfix10_En0 
 input [9:0] Pix_270, // sfix10_En0 
 input [9:0] Pix_271, // sfix10_En0 
 input [9:0] Pix_272, // sfix10_En0 
 input [9:0] Pix_273, // sfix10_En0 
 input [9:0] Pix_274, // sfix10_En0 
 input [9:0] Pix_275, // sfix10_En0 
 input [9:0] Pix_276, // sfix10_En0 
 input [9:0] Pix_277, // sfix10_En0 
 input [9:0] Pix_278, // sfix10_En0 
 input [9:0] Pix_279, // sfix10_En0 
 input [9:0] Pix_280, // sfix10_En0 
 input [9:0] Pix_281, // sfix10_En0 
 input [9:0] Pix_282, // sfix10_En0 
 input [9:0] Pix_283, // sfix10_En0 
 input [9:0] Pix_284, // sfix10_En0 
 input [9:0] Pix_285, // sfix10_En0 
 input [9:0] Pix_286, // sfix10_En0 
 input [9:0] Pix_287, // sfix10_En0 
 input [9:0] Pix_288, // sfix10_En0 
 input [9:0] Pix_289, // sfix10_En0 
 input [9:0] Pix_290, // sfix10_En0 
 input [9:0] Pix_291, // sfix10_En0 
 input [9:0] Pix_292, // sfix10_En0 
 input [9:0] Pix_293, // sfix10_En0 
 input [9:0] Pix_294, // sfix10_En0 
 input [9:0] Pix_295, // sfix10_En0 
 input [9:0] Pix_296, // sfix10_En0 
 input [9:0] Pix_297, // sfix10_En0 
 input [9:0] Pix_298, // sfix10_En0 
 input [9:0] Pix_299, // sfix10_En0 
 input [9:0] Pix_300, // sfix10_En0 
 input [9:0] Pix_301, // sfix10_En0 
 input [9:0] Pix_302, // sfix10_En0 
 input [9:0] Pix_303, // sfix10_En0 
 input [9:0] Pix_304, // sfix10_En0 
 input [9:0] Pix_305, // sfix10_En0 
 input [9:0] Pix_306, // sfix10_En0 
 input [9:0] Pix_307, // sfix10_En0 
 input [9:0] Pix_308, // sfix10_En0 
 input [9:0] Pix_309, // sfix10_En0 
 input [9:0] Pix_310, // sfix10_En0 
 input [9:0] Pix_311, // sfix10_En0 
 input [9:0] Pix_312, // sfix10_En0 
 input [9:0] Pix_313, // sfix10_En0 
 input [9:0] Pix_314, // sfix10_En0 
 input [9:0] Pix_315, // sfix10_En0 
 input [9:0] Pix_316, // sfix10_En0 
 input [9:0] Pix_317, // sfix10_En0 
 input [9:0] Pix_318, // sfix10_En0 
 input [9:0] Pix_319, // sfix10_En0 
 input [9:0] Pix_320, // sfix10_En0 
 input [9:0] Pix_321, // sfix10_En0 
 input [9:0] Pix_322, // sfix10_En0 
 input [9:0] Pix_323, // sfix10_En0 
 input [9:0] Pix_324, // sfix10_En0 
 input [9:0] Pix_325, // sfix10_En0 
 input [9:0] Pix_326, // sfix10_En0 
 input [9:0] Pix_327, // sfix10_En0 
 input [9:0] Pix_328, // sfix10_En0 
 input [9:0] Pix_329, // sfix10_En0 
 input [9:0] Pix_330, // sfix10_En0 
 input [9:0] Pix_331, // sfix10_En0 
 input [9:0] Pix_332, // sfix10_En0 
 input [9:0] Pix_333, // sfix10_En0 
 input [9:0] Pix_334, // sfix10_En0 
 input [9:0] Pix_335, // sfix10_En0 
 input [9:0] Pix_336, // sfix10_En0 
 input [9:0] Pix_337, // sfix10_En0 
 input [9:0] Pix_338, // sfix10_En0 
 input [9:0] Pix_339, // sfix10_En0 
 input [9:0] Pix_340, // sfix10_En0 
 input [9:0] Pix_341, // sfix10_En0 
 input [9:0] Pix_342, // sfix10_En0 
 input [9:0] Pix_343, // sfix10_En0 
 input [9:0] Pix_344, // sfix10_En0 
 input [9:0] Pix_345, // sfix10_En0 
 input [9:0] Pix_346, // sfix10_En0 
 input [9:0] Pix_347, // sfix10_En0 
 input [9:0] Pix_348, // sfix10_En0 
 input [9:0] Pix_349, // sfix10_En0 
 input [9:0] Pix_350, // sfix10_En0 
 input [9:0] Pix_351, // sfix10_En0 
 input [9:0] Pix_352, // sfix10_En0 
 input [9:0] Pix_353, // sfix10_En0 
 input [9:0] Pix_354, // sfix10_En0 
 input [9:0] Pix_355, // sfix10_En0 
 input [9:0] Pix_356, // sfix10_En0 
 input [9:0] Pix_357, // sfix10_En0 
 input [9:0] Pix_358, // sfix10_En0 
 input [9:0] Pix_359, // sfix10_En0 
 input [9:0] Pix_360, // sfix10_En0 
 input [9:0] Pix_361, // sfix10_En0 
 input [9:0] Pix_362, // sfix10_En0 
 input [9:0] Pix_363, // sfix10_En0 
 input [9:0] Pix_364, // sfix10_En0 
 input [9:0] Pix_365, // sfix10_En0 
 input [9:0] Pix_366, // sfix10_En0 
 input [9:0] Pix_367, // sfix10_En0 
 input [9:0] Pix_368, // sfix10_En0 
 input [9:0] Pix_369, // sfix10_En0 
 input [9:0] Pix_370, // sfix10_En0 
 input [9:0] Pix_371, // sfix10_En0 
 input [9:0] Pix_372, // sfix10_En0 
 input [9:0] Pix_373, // sfix10_En0 
 input [9:0] Pix_374, // sfix10_En0 
 input [9:0] Pix_375, // sfix10_En0 
 input [9:0] Pix_376, // sfix10_En0 
 input [9:0] Pix_377, // sfix10_En0 
 input [9:0] Pix_378, // sfix10_En0 
 input [9:0] Pix_379, // sfix10_En0 
 input [9:0] Pix_380, // sfix10_En0 
 input [9:0] Pix_381, // sfix10_En0 
 input [9:0] Pix_382, // sfix10_En0 
 input [9:0] Pix_383, // sfix10_En0 
 input [9:0] Pix_384, // sfix10_En0 
 input [9:0] Pix_385, // sfix10_En0 
 input [9:0] Pix_386, // sfix10_En0 
 input [9:0] Pix_387, // sfix10_En0 
 input [9:0] Pix_388, // sfix10_En0 
 input [9:0] Pix_389, // sfix10_En0 
 input [9:0] Pix_390, // sfix10_En0 
 input [9:0] Pix_391, // sfix10_En0 
 input [9:0] Pix_392, // sfix10_En0 
 input [9:0] Pix_393, // sfix10_En0 
 input [9:0] Pix_394, // sfix10_En0 
 input [9:0] Pix_395, // sfix10_En0 
 input [9:0] Pix_396, // sfix10_En0 
 input [9:0] Pix_397, // sfix10_En0 
 input [9:0] Pix_398, // sfix10_En0 
 input [9:0] Pix_399, // sfix10_En0 
 input [9:0] Pix_400, // sfix10_En0 
 input [9:0] Pix_401, // sfix10_En0 
 input [9:0] Pix_402, // sfix10_En0 
 input [9:0] Pix_403, // sfix10_En0 
 input [9:0] Pix_404, // sfix10_En0 
 input [9:0] Pix_405, // sfix10_En0 
 input [9:0] Pix_406, // sfix10_En0 
 input [9:0] Pix_407, // sfix10_En0 
 input [9:0] Pix_408, // sfix10_En0 
 input [9:0] Pix_409, // sfix10_En0 
 input [9:0] Pix_410, // sfix10_En0 
 input [9:0] Pix_411, // sfix10_En0 
 input [9:0] Pix_412, // sfix10_En0 
 input [9:0] Pix_413, // sfix10_En0 
 input [9:0] Pix_414, // sfix10_En0 
 input [9:0] Pix_415, // sfix10_En0 
 input [9:0] Pix_416, // sfix10_En0 
 input [9:0] Pix_417, // sfix10_En0 
 input [9:0] Pix_418, // sfix10_En0 
 input [9:0] Pix_419, // sfix10_En0 
 input [9:0] Pix_420, // sfix10_En0 
 input [9:0] Pix_421, // sfix10_En0 
 input [9:0] Pix_422, // sfix10_En0 
 input [9:0] Pix_423, // sfix10_En0 
 input [9:0] Pix_424, // sfix10_En0 
 input [9:0] Pix_425, // sfix10_En0 
 input [9:0] Pix_426, // sfix10_En0 
 input [9:0] Pix_427, // sfix10_En0 
 input [9:0] Pix_428, // sfix10_En0 
 input [9:0] Pix_429, // sfix10_En0 
 input [9:0] Pix_430, // sfix10_En0 
 input [9:0] Pix_431, // sfix10_En0 
 input [9:0] Pix_432, // sfix10_En0 
 input [9:0] Pix_433, // sfix10_En0 
 input [9:0] Pix_434, // sfix10_En0 
 input [9:0] Pix_435, // sfix10_En0 
 input [9:0] Pix_436, // sfix10_En0 
 input [9:0] Pix_437, // sfix10_En0 
 input [9:0] Pix_438, // sfix10_En0 
 input [9:0] Pix_439, // sfix10_En0 
 input [9:0] Pix_440, // sfix10_En0 
 input [9:0] Pix_441, // sfix10_En0 
 input [9:0] Pix_442, // sfix10_En0 
 input [9:0] Pix_443, // sfix10_En0 
 input [9:0] Pix_444, // sfix10_En0 
 input [9:0] Pix_445, // sfix10_En0 
 input [9:0] Pix_446, // sfix10_En0 
 input [9:0] Pix_447, // sfix10_En0 
 input [9:0] Pix_448, // sfix10_En0 
 input [9:0] Pix_449, // sfix10_En0 
 input [9:0] Pix_450, // sfix10_En0 
 input [9:0] Pix_451, // sfix10_En0 
 input [9:0] Pix_452, // sfix10_En0 
 input [9:0] Pix_453, // sfix10_En0 
 input [9:0] Pix_454, // sfix10_En0 
 input [9:0] Pix_455, // sfix10_En0 
 input [9:0] Pix_456, // sfix10_En0 
 input [9:0] Pix_457, // sfix10_En0 
 input [9:0] Pix_458, // sfix10_En0 
 input [9:0] Pix_459, // sfix10_En0 
 input [9:0] Pix_460, // sfix10_En0 
 input [9:0] Pix_461, // sfix10_En0 
 input [9:0] Pix_462, // sfix10_En0 
 input [9:0] Pix_463, // sfix10_En0 
 input [9:0] Pix_464, // sfix10_En0 
 input [9:0] Pix_465, // sfix10_En0 
 input [9:0] Pix_466, // sfix10_En0 
 input [9:0] Pix_467, // sfix10_En0 
 input [9:0] Pix_468, // sfix10_En0 
 input [9:0] Pix_469, // sfix10_En0 
 input [9:0] Pix_470, // sfix10_En0 
 input [9:0] Pix_471, // sfix10_En0 
 input [9:0] Pix_472, // sfix10_En0 
 input [9:0] Pix_473, // sfix10_En0 
 input [9:0] Pix_474, // sfix10_En0 
 input [9:0] Pix_475, // sfix10_En0 
 input [9:0] Pix_476, // sfix10_En0 
 input [9:0] Pix_477, // sfix10_En0 
 input [9:0] Pix_478, // sfix10_En0 
 input [9:0] Pix_479, // sfix10_En0 
 input [9:0] Pix_480, // sfix10_En0 
 input [9:0] Pix_481, // sfix10_En0 
 input [9:0] Pix_482, // sfix10_En0 
 input [9:0] Pix_483, // sfix10_En0 
 input [9:0] Pix_484, // sfix10_En0 
 input [9:0] Pix_485, // sfix10_En0 
 input [9:0] Pix_486, // sfix10_En0 
 input [9:0] Pix_487, // sfix10_En0 
 input [9:0] Pix_488, // sfix10_En0 
 input [9:0] Pix_489, // sfix10_En0 
 input [9:0] Pix_490, // sfix10_En0 
 input [9:0] Pix_491, // sfix10_En0 
 input [9:0] Pix_492, // sfix10_En0 
 input [9:0] Pix_493, // sfix10_En0 
 input [9:0] Pix_494, // sfix10_En0 
 input [9:0] Pix_495, // sfix10_En0 
 input [9:0] Pix_496, // sfix10_En0 
 input [9:0] Pix_497, // sfix10_En0 
 input [9:0] Pix_498, // sfix10_En0 
 input [9:0] Pix_499, // sfix10_En0 
 input [9:0] Pix_500, // sfix10_En0 
 input [9:0] Pix_501, // sfix10_En0 
 input [9:0] Pix_502, // sfix10_En0 
 input [9:0] Pix_503, // sfix10_En0 
 input [9:0] Pix_504, // sfix10_En0 
 input [9:0] Pix_505, // sfix10_En0 
 input [9:0] Pix_506, // sfix10_En0 
 input [9:0] Pix_507, // sfix10_En0 
 input [9:0] Pix_508, // sfix10_En0 
 input [9:0] Pix_509, // sfix10_En0 
 input [9:0] Pix_510, // sfix10_En0 
 input [9:0] Pix_511, // sfix10_En0 
 input [9:0] Pix_512, // sfix10_En0 
 input [9:0] Pix_513, // sfix10_En0 
 input [9:0] Pix_514, // sfix10_En0 
 input [9:0] Pix_515, // sfix10_En0 
 input [9:0] Pix_516, // sfix10_En0 
 input [9:0] Pix_517, // sfix10_En0 
 input [9:0] Pix_518, // sfix10_En0 
 input [9:0] Pix_519, // sfix10_En0 
 input [9:0] Pix_520, // sfix10_En0 
 input [9:0] Pix_521, // sfix10_En0 
 input [9:0] Pix_522, // sfix10_En0 
 input [9:0] Pix_523, // sfix10_En0 
 input [9:0] Pix_524, // sfix10_En0 
 input [9:0] Pix_525, // sfix10_En0 
 input [9:0] Pix_526, // sfix10_En0 
 input [9:0] Pix_527, // sfix10_En0 
 input [9:0] Pix_528, // sfix10_En0 
 input [9:0] Pix_529, // sfix10_En0 
 input [9:0] Pix_530, // sfix10_En0 
 input [9:0] Pix_531, // sfix10_En0 
 input [9:0] Pix_532, // sfix10_En0 
 input [9:0] Pix_533, // sfix10_En0 
 input [9:0] Pix_534, // sfix10_En0 
 input [9:0] Pix_535, // sfix10_En0 
 input [9:0] Pix_536, // sfix10_En0 
 input [9:0] Pix_537, // sfix10_En0 
 input [9:0] Pix_538, // sfix10_En0 
 input [9:0] Pix_539, // sfix10_En0 
 input [9:0] Pix_540, // sfix10_En0 
 input [9:0] Pix_541, // sfix10_En0 
 input [9:0] Pix_542, // sfix10_En0 
 input [9:0] Pix_543, // sfix10_En0 
 input [9:0] Pix_544, // sfix10_En0 
 input [9:0] Pix_545, // sfix10_En0 
 input [9:0] Pix_546, // sfix10_En0 
 input [9:0] Pix_547, // sfix10_En0 
 input [9:0] Pix_548, // sfix10_En0 
 input [9:0] Pix_549, // sfix10_En0 
 input [9:0] Pix_550, // sfix10_En0 
 input [9:0] Pix_551, // sfix10_En0 
 input [9:0] Pix_552, // sfix10_En0 
 input [9:0] Pix_553, // sfix10_En0 
 input [9:0] Pix_554, // sfix10_En0 
 input [9:0] Pix_555, // sfix10_En0 
 input [9:0] Pix_556, // sfix10_En0 
 input [9:0] Pix_557, // sfix10_En0 
 input [9:0] Pix_558, // sfix10_En0 
 input [9:0] Pix_559, // sfix10_En0 
 input [9:0] Pix_560, // sfix10_En0 
 input [9:0] Pix_561, // sfix10_En0 
 input [9:0] Pix_562, // sfix10_En0 
 input [9:0] Pix_563, // sfix10_En0 
 input [9:0] Pix_564, // sfix10_En0 
 input [9:0] Pix_565, // sfix10_En0 
 input [9:0] Pix_566, // sfix10_En0 
 input [9:0] Pix_567, // sfix10_En0 
 input [9:0] Pix_568, // sfix10_En0 
 input [9:0] Pix_569, // sfix10_En0 
 input [9:0] Pix_570, // sfix10_En0 
 input [9:0] Pix_571, // sfix10_En0 
 input [9:0] Pix_572, // sfix10_En0 
 input [9:0] Pix_573, // sfix10_En0 
 input [9:0] Pix_574, // sfix10_En0 
 input [9:0] Pix_575, // sfix10_En0 
 input [9:0] Pix_576, // sfix10_En0 
 input [9:0] Pix_577, // sfix10_En0 
 input [9:0] Pix_578, // sfix10_En0 
 input [9:0] Pix_579, // sfix10_En0 
 input [9:0] Pix_580, // sfix10_En0 
 input [9:0] Pix_581, // sfix10_En0 
 input [9:0] Pix_582, // sfix10_En0 
 input [9:0] Pix_583, // sfix10_En0 
 input [9:0] Pix_584, // sfix10_En0 
 input [9:0] Pix_585, // sfix10_En0 
 input [9:0] Pix_586, // sfix10_En0 
 input [9:0] Pix_587, // sfix10_En0 
 input [9:0] Pix_588, // sfix10_En0 
 input [9:0] Pix_589, // sfix10_En0 
 input [9:0] Pix_590, // sfix10_En0 
 input [9:0] Pix_591, // sfix10_En0 
 input [9:0] Pix_592, // sfix10_En0 
 input [9:0] Pix_593, // sfix10_En0 
 input [9:0] Pix_594, // sfix10_En0 
 input [9:0] Pix_595, // sfix10_En0 
 input [9:0] Pix_596, // sfix10_En0 
 input [9:0] Pix_597, // sfix10_En0 
 input [9:0] Pix_598, // sfix10_En0 
 input [9:0] Pix_599, // sfix10_En0 
 input [9:0] Pix_600, // sfix10_En0 
 input [9:0] Pix_601, // sfix10_En0 
 input [9:0] Pix_602, // sfix10_En0 
 input [9:0] Pix_603, // sfix10_En0 
 input [9:0] Pix_604, // sfix10_En0 
 input [9:0] Pix_605, // sfix10_En0 
 input [9:0] Pix_606, // sfix10_En0 
 input [9:0] Pix_607, // sfix10_En0 
 input [9:0] Pix_608, // sfix10_En0 
 input [9:0] Pix_609, // sfix10_En0 
 input [9:0] Pix_610, // sfix10_En0 
 input [9:0] Pix_611, // sfix10_En0 
 input [9:0] Pix_612, // sfix10_En0 
 input [9:0] Pix_613, // sfix10_En0 
 input [9:0] Pix_614, // sfix10_En0 
 input [9:0] Pix_615, // sfix10_En0 
 input [9:0] Pix_616, // sfix10_En0 
 input [9:0] Pix_617, // sfix10_En0 
 input [9:0] Pix_618, // sfix10_En0 
 input [9:0] Pix_619, // sfix10_En0 
 input [9:0] Pix_620, // sfix10_En0 
 input [9:0] Pix_621, // sfix10_En0 
 input [9:0] Pix_622, // sfix10_En0 
 input [9:0] Pix_623, // sfix10_En0 
 input [9:0] Pix_624, // sfix10_En0 
 input [9:0] Pix_625, // sfix10_En0 
 input [9:0] Pix_626, // sfix10_En0 
 input [9:0] Pix_627, // sfix10_En0 
 input [9:0] Pix_628, // sfix10_En0 
 input [9:0] Pix_629, // sfix10_En0 
 input [9:0] Pix_630, // sfix10_En0 
 input [9:0] Pix_631, // sfix10_En0 
 input [9:0] Pix_632, // sfix10_En0 
 input [9:0] Pix_633, // sfix10_En0 
 input [9:0] Pix_634, // sfix10_En0 
 input [9:0] Pix_635, // sfix10_En0 
 input [9:0] Pix_636, // sfix10_En0 
 input [9:0] Pix_637, // sfix10_En0 
 input [9:0] Pix_638, // sfix10_En0 
 input [9:0] Pix_639, // sfix10_En0 
 input [9:0] Pix_640, // sfix10_En0 
 input [9:0] Pix_641, // sfix10_En0 
 input [9:0] Pix_642, // sfix10_En0 
 input [9:0] Pix_643, // sfix10_En0 
 input [9:0] Pix_644, // sfix10_En0 
 input [9:0] Pix_645, // sfix10_En0 
 input [9:0] Pix_646, // sfix10_En0 
 input [9:0] Pix_647, // sfix10_En0 
 input [9:0] Pix_648, // sfix10_En0 
 input [9:0] Pix_649, // sfix10_En0 
 input [9:0] Pix_650, // sfix10_En0 
 input [9:0] Pix_651, // sfix10_En0 
 input [9:0] Pix_652, // sfix10_En0 
 input [9:0] Pix_653, // sfix10_En0 
 input [9:0] Pix_654, // sfix10_En0 
 input [9:0] Pix_655, // sfix10_En0 
 input [9:0] Pix_656, // sfix10_En0 
 input [9:0] Pix_657, // sfix10_En0 
 input [9:0] Pix_658, // sfix10_En0 
 input [9:0] Pix_659, // sfix10_En0 
 input [9:0] Pix_660, // sfix10_En0 
 input [9:0] Pix_661, // sfix10_En0 
 input [9:0] Pix_662, // sfix10_En0 
 input [9:0] Pix_663, // sfix10_En0 
 input [9:0] Pix_664, // sfix10_En0 
 input [9:0] Pix_665, // sfix10_En0 
 input [9:0] Pix_666, // sfix10_En0 
 input [9:0] Pix_667, // sfix10_En0 
 input [9:0] Pix_668, // sfix10_En0 
 input [9:0] Pix_669, // sfix10_En0 
 input [9:0] Pix_670, // sfix10_En0 
 input [9:0] Pix_671, // sfix10_En0 
 input [9:0] Pix_672, // sfix10_En0 
 input [9:0] Pix_673, // sfix10_En0 
 input [9:0] Pix_674, // sfix10_En0 
 input [9:0] Pix_675, // sfix10_En0 
 input [9:0] Pix_676, // sfix10_En0 
 input [9:0] Pix_677, // sfix10_En0 
 input [9:0] Pix_678, // sfix10_En0 
 input [9:0] Pix_679, // sfix10_En0 
 input [9:0] Pix_680, // sfix10_En0 
 input [9:0] Pix_681, // sfix10_En0 
 input [9:0] Pix_682, // sfix10_En0 
 input [9:0] Pix_683, // sfix10_En0 
 input [9:0] Pix_684, // sfix10_En0 
 input [9:0] Pix_685, // sfix10_En0 
 input [9:0] Pix_686, // sfix10_En0 
 input [9:0] Pix_687, // sfix10_En0 
 input [9:0] Pix_688, // sfix10_En0 
 input [9:0] Pix_689, // sfix10_En0 
 input [9:0] Pix_690, // sfix10_En0 
 input [9:0] Pix_691, // sfix10_En0 
 input [9:0] Pix_692, // sfix10_En0 
 input [9:0] Pix_693, // sfix10_En0 
 input [9:0] Pix_694, // sfix10_En0 
 input [9:0] Pix_695, // sfix10_En0 
 input [9:0] Pix_696, // sfix10_En0 
 input [9:0] Pix_697, // sfix10_En0 
 input [9:0] Pix_698, // sfix10_En0 
 input [9:0] Pix_699, // sfix10_En0 
 input [9:0] Pix_700, // sfix10_En0 
 input [9:0] Pix_701, // sfix10_En0 
 input [9:0] Pix_702, // sfix10_En0 
 input [9:0] Pix_703, // sfix10_En0 
 input [9:0] Pix_704, // sfix10_En0 
 input [9:0] Pix_705, // sfix10_En0 
 input [9:0] Pix_706, // sfix10_En0 
 input [9:0] Pix_707, // sfix10_En0 
 input [9:0] Pix_708, // sfix10_En0 
 input [9:0] Pix_709, // sfix10_En0 
 input [9:0] Pix_710, // sfix10_En0 
 input [9:0] Pix_711, // sfix10_En0 
 input [9:0] Pix_712, // sfix10_En0 
 input [9:0] Pix_713, // sfix10_En0 
 input [9:0] Pix_714, // sfix10_En0 
 input [9:0] Pix_715, // sfix10_En0 
 input [9:0] Pix_716, // sfix10_En0 
 input [9:0] Pix_717, // sfix10_En0 
 input [9:0] Pix_718, // sfix10_En0 
 input [9:0] Pix_719, // sfix10_En0 
 input [9:0] Pix_720, // sfix10_En0 
 input [9:0] Pix_721, // sfix10_En0 
 input [9:0] Pix_722, // sfix10_En0 
 input [9:0] Pix_723, // sfix10_En0 
 input [9:0] Pix_724, // sfix10_En0 
 input [9:0] Pix_725, // sfix10_En0 
 input [9:0] Pix_726, // sfix10_En0 
 input [9:0] Pix_727, // sfix10_En0 
 input [9:0] Pix_728, // sfix10_En0 
 input [9:0] Pix_729, // sfix10_En0 
 input [9:0] Pix_730, // sfix10_En0 
 input [9:0] Pix_731, // sfix10_En0 
 input [9:0] Pix_732, // sfix10_En0 
 input [9:0] Pix_733, // sfix10_En0 
 input [9:0] Pix_734, // sfix10_En0 
 input [9:0] Pix_735, // sfix10_En0 
 input [9:0] Pix_736, // sfix10_En0 
 input [9:0] Pix_737, // sfix10_En0 
 input [9:0] Pix_738, // sfix10_En0 
 input [9:0] Pix_739, // sfix10_En0 
 input [9:0] Pix_740, // sfix10_En0 
 input [9:0] Pix_741, // sfix10_En0 
 input [9:0] Pix_742, // sfix10_En0 
 input [9:0] Pix_743, // sfix10_En0 
 input [9:0] Pix_744, // sfix10_En0 
 input [9:0] Pix_745, // sfix10_En0 
 input [9:0] Pix_746, // sfix10_En0 
 input [9:0] Pix_747, // sfix10_En0 
 input [9:0] Pix_748, // sfix10_En0 
 input [9:0] Pix_749, // sfix10_En0 
 input [9:0] Pix_750, // sfix10_En0 
 input [9:0] Pix_751, // sfix10_En0 
 input [9:0] Pix_752, // sfix10_En0 
 input [9:0] Pix_753, // sfix10_En0 
 input [9:0] Pix_754, // sfix10_En0 
 input [9:0] Pix_755, // sfix10_En0 
 input [9:0] Pix_756, // sfix10_En0 
 input [9:0] Pix_757, // sfix10_En0 
 input [9:0] Pix_758, // sfix10_En0 
 input [9:0] Pix_759, // sfix10_En0 
 input [9:0] Pix_760, // sfix10_En0 
 input [9:0] Pix_761, // sfix10_En0 
 input [9:0] Pix_762, // sfix10_En0 
 input [9:0] Pix_763, // sfix10_En0 
 input [9:0] Pix_764, // sfix10_En0 
 input [9:0] Pix_765, // sfix10_En0 
 input [9:0] Pix_766, // sfix10_En0 
 input [9:0] Pix_767, // sfix10_En0 
 input [9:0] Pix_768, // sfix10_En0 
 input [9:0] Pix_769, // sfix10_En0 
 input [9:0] Pix_770, // sfix10_En0 
 input [9:0] Pix_771, // sfix10_En0 
 input [9:0] Pix_772, // sfix10_En0 
 input [9:0] Pix_773, // sfix10_En0 
 input [9:0] Pix_774, // sfix10_En0 
 input [9:0] Pix_775, // sfix10_En0 
 input [9:0] Pix_776, // sfix10_En0 
 input [9:0] Pix_777, // sfix10_En0 
 input [9:0] Pix_778, // sfix10_En0 
 input [9:0] Pix_779, // sfix10_En0 
 input [9:0] Pix_780, // sfix10_En0 
 input [9:0] Pix_781, // sfix10_En0 
 input [9:0] Pix_782, // sfix10_En0 
 input [9:0] Pix_783, // sfix10_En0 
 input [9:0] Pix_784, // sfix10_En0 
 output [3:0] Image_Number, // sfix26_En18 
 output Output_Valid 
);

//--------------------------------------------------------------------------------------------------------------------------------------------------
//input register
reg [18:0] w_0_0,w_0_1,w_0_2,w_0_3,w_0_4,w_0_5,w_0_6,w_0_7,w_0_8,w_0_9,w_0_10,w_0_11,w_0_12,w_0_13,w_0_14,w_0_15,w_0_16,w_0_17,w_0_18,w_0_19,w_0_20,w_0_21,w_0_22,w_0_23,w_0_24,w_0_25,w_0_26,w_0_27,w_0_28,w_0_29,w_0_30,w_0_31,w_0_32,w_0_33,w_0_34,w_0_35,w_0_36,w_0_37,w_0_38,w_0_39,w_0_40,w_0_41,w_0_42,w_0_43,w_0_44,w_0_45,w_0_46,w_0_47,w_0_48,w_0_49,w_0_50,w_0_51,w_0_52,w_0_53,w_0_54,w_0_55,w_0_56,w_0_57,w_0_58,w_0_59,w_0_60,w_0_61,w_0_62,w_0_63,w_0_64,w_0_65,w_0_66,w_0_67,w_0_68,w_0_69,w_0_70,w_0_71,w_0_72,w_0_73,w_0_74,w_0_75,w_0_76,w_0_77,w_0_78,w_0_79,w_0_80,w_0_81,w_0_82,w_0_83,w_0_84,w_0_85,w_0_86,w_0_87,w_0_88,w_0_89,w_0_90,w_0_91,w_0_92,w_0_93,w_0_94,w_0_95,w_0_96,w_0_97,w_0_98,w_0_99,w_0_100,w_0_101,w_0_102,w_0_103,w_0_104,w_0_105,w_0_106,w_0_107,w_0_108,w_0_109,w_0_110,w_0_111,w_0_112,w_0_113,w_0_114,w_0_115,w_0_116,w_0_117,w_0_118,w_0_119,w_0_120,w_0_121,w_0_122,w_0_123,w_0_124,w_0_125,w_0_126,w_0_127,w_0_128,w_0_129,w_0_130,w_0_131,w_0_132,w_0_133,w_0_134,w_0_135,w_0_136,w_0_137,w_0_138,w_0_139,w_0_140,w_0_141,w_0_142,w_0_143,w_0_144,w_0_145,w_0_146,w_0_147,w_0_148,w_0_149,w_0_150,w_0_151,w_0_152,w_0_153,w_0_154,w_0_155,w_0_156,w_0_157,w_0_158,w_0_159,w_0_160,w_0_161,w_0_162,w_0_163,w_0_164,w_0_165,w_0_166,w_0_167,w_0_168,w_0_169,w_0_170,w_0_171,w_0_172,w_0_173,w_0_174,w_0_175,w_0_176,w_0_177,w_0_178,w_0_179,w_0_180,w_0_181,w_0_182,w_0_183,w_0_184,w_0_185,w_0_186,w_0_187,w_0_188,w_0_189,w_0_190,w_0_191,w_0_192,w_0_193,w_0_194,w_0_195,w_0_196,w_0_197,w_0_198,w_0_199,w_0_200,w_0_201,w_0_202,w_0_203,w_0_204,w_0_205,w_0_206,w_0_207,w_0_208,w_0_209,w_0_210,w_0_211,w_0_212,w_0_213,w_0_214,w_0_215,w_0_216,w_0_217,w_0_218,w_0_219,w_0_220,w_0_221,w_0_222,w_0_223,w_0_224,w_0_225,w_0_226,w_0_227,w_0_228,w_0_229,w_0_230,w_0_231,w_0_232,w_0_233,w_0_234,w_0_235,w_0_236,w_0_237,w_0_238,w_0_239,w_0_240,w_0_241,w_0_242,w_0_243,w_0_244,w_0_245,w_0_246,w_0_247,w_0_248,w_0_249,w_0_250,w_0_251,w_0_252,w_0_253,w_0_254,w_0_255,w_0_256,w_0_257,w_0_258,w_0_259,w_0_260,w_0_261,w_0_262,w_0_263,w_0_264,w_0_265,w_0_266,w_0_267,w_0_268,w_0_269,w_0_270,w_0_271,w_0_272,w_0_273,w_0_274,w_0_275,w_0_276,w_0_277,w_0_278,w_0_279,w_0_280,w_0_281,w_0_282,w_0_283,w_0_284,w_0_285,w_0_286,w_0_287,w_0_288,w_0_289,w_0_290,w_0_291,w_0_292,w_0_293,w_0_294,w_0_295,w_0_296,w_0_297,w_0_298,w_0_299,w_0_300,w_0_301,w_0_302,w_0_303,w_0_304,w_0_305,w_0_306,w_0_307,w_0_308,w_0_309,w_0_310,w_0_311,w_0_312,w_0_313,w_0_314,w_0_315,w_0_316,w_0_317,w_0_318,w_0_319,w_0_320,w_0_321,w_0_322,w_0_323,w_0_324,w_0_325,w_0_326,w_0_327,w_0_328,w_0_329,w_0_330,w_0_331,w_0_332,w_0_333,w_0_334,w_0_335,w_0_336,w_0_337,w_0_338,w_0_339,w_0_340,w_0_341,w_0_342,w_0_343,w_0_344,w_0_345,w_0_346,w_0_347,w_0_348,w_0_349,w_0_350,w_0_351,w_0_352,w_0_353,w_0_354,w_0_355,w_0_356,w_0_357,w_0_358,w_0_359,w_0_360,w_0_361,w_0_362,w_0_363,w_0_364,w_0_365,w_0_366,w_0_367,w_0_368,w_0_369,w_0_370,w_0_371,w_0_372,w_0_373,w_0_374,w_0_375,w_0_376,w_0_377,w_0_378,w_0_379,w_0_380,w_0_381,w_0_382,w_0_383,w_0_384,w_0_385,w_0_386,w_0_387,w_0_388,w_0_389,w_0_390,w_0_391,w_0_392,w_0_393,w_0_394,w_0_395,w_0_396,w_0_397,w_0_398,w_0_399,w_0_400,w_0_401,w_0_402,w_0_403,w_0_404,w_0_405,w_0_406,w_0_407,w_0_408,w_0_409,w_0_410,w_0_411,w_0_412,w_0_413,w_0_414,w_0_415,w_0_416,w_0_417,w_0_418,w_0_419,w_0_420,w_0_421,w_0_422,w_0_423,w_0_424,w_0_425,w_0_426,w_0_427,w_0_428,w_0_429,w_0_430,w_0_431,w_0_432,w_0_433,w_0_434,w_0_435,w_0_436,w_0_437,w_0_438,w_0_439,w_0_440,w_0_441,w_0_442,w_0_443,w_0_444,w_0_445,w_0_446,w_0_447,w_0_448,w_0_449,w_0_450,w_0_451,w_0_452,w_0_453,w_0_454,w_0_455,w_0_456,w_0_457,w_0_458,w_0_459,w_0_460,w_0_461,w_0_462,w_0_463,w_0_464,w_0_465,w_0_466,w_0_467,w_0_468,w_0_469,w_0_470,w_0_471,w_0_472,w_0_473,w_0_474,w_0_475,w_0_476,w_0_477,w_0_478,w_0_479,w_0_480,w_0_481,w_0_482,w_0_483,w_0_484,w_0_485,w_0_486,w_0_487,w_0_488,w_0_489,w_0_490,w_0_491,w_0_492,w_0_493,w_0_494,w_0_495,w_0_496,w_0_497,w_0_498,w_0_499,w_0_500,w_0_501,w_0_502,w_0_503,w_0_504,w_0_505,w_0_506,w_0_507,w_0_508,w_0_509,w_0_510,w_0_511,w_0_512,w_0_513,w_0_514,w_0_515,w_0_516,w_0_517,w_0_518,w_0_519,w_0_520,w_0_521,w_0_522,w_0_523,w_0_524,w_0_525,w_0_526,w_0_527,w_0_528,w_0_529,w_0_530,w_0_531,w_0_532,w_0_533,w_0_534,w_0_535,w_0_536,w_0_537,w_0_538,w_0_539,w_0_540,w_0_541,w_0_542,w_0_543,w_0_544,w_0_545,w_0_546,w_0_547,w_0_548,w_0_549,w_0_550,w_0_551,w_0_552,w_0_553,w_0_554,w_0_555,w_0_556,w_0_557,w_0_558,w_0_559,w_0_560,w_0_561,w_0_562,w_0_563,w_0_564,w_0_565,w_0_566,w_0_567,w_0_568,w_0_569,w_0_570,w_0_571,w_0_572,w_0_573,w_0_574,w_0_575,w_0_576,w_0_577,w_0_578,w_0_579,w_0_580,w_0_581,w_0_582,w_0_583,w_0_584,w_0_585,w_0_586,w_0_587,w_0_588,w_0_589,w_0_590,w_0_591,w_0_592,w_0_593,w_0_594,w_0_595,w_0_596,w_0_597,w_0_598,w_0_599,w_0_600,w_0_601,w_0_602,w_0_603,w_0_604,w_0_605,w_0_606,w_0_607,w_0_608,w_0_609,w_0_610,w_0_611,w_0_612,w_0_613,w_0_614,w_0_615,w_0_616,w_0_617,w_0_618,w_0_619,w_0_620,w_0_621,w_0_622,w_0_623,w_0_624,w_0_625,w_0_626,w_0_627,w_0_628,w_0_629,w_0_630,w_0_631,w_0_632,w_0_633,w_0_634,w_0_635,w_0_636,w_0_637,w_0_638,w_0_639,w_0_640,w_0_641,w_0_642,w_0_643,w_0_644,w_0_645,w_0_646,w_0_647,w_0_648,w_0_649,w_0_650,w_0_651,w_0_652,w_0_653,w_0_654,w_0_655,w_0_656,w_0_657,w_0_658,w_0_659,w_0_660,w_0_661,w_0_662,w_0_663,w_0_664,w_0_665,w_0_666,w_0_667,w_0_668,w_0_669,w_0_670,w_0_671,w_0_672,w_0_673,w_0_674,w_0_675,w_0_676,w_0_677,w_0_678,w_0_679,w_0_680,w_0_681,w_0_682,w_0_683,w_0_684,w_0_685,w_0_686,w_0_687,w_0_688,w_0_689,w_0_690,w_0_691,w_0_692,w_0_693,w_0_694,w_0_695,w_0_696,w_0_697,w_0_698,w_0_699,w_0_700,w_0_701,w_0_702,w_0_703,w_0_704,w_0_705,w_0_706,w_0_707,w_0_708,w_0_709,w_0_710,w_0_711,w_0_712,w_0_713,w_0_714,w_0_715,w_0_716,w_0_717,w_0_718,w_0_719,w_0_720,w_0_721,w_0_722,w_0_723,w_0_724,w_0_725,w_0_726,w_0_727,w_0_728,w_0_729,w_0_730,w_0_731,w_0_732,w_0_733,w_0_734,w_0_735,w_0_736,w_0_737,w_0_738,w_0_739,w_0_740,w_0_741,w_0_742,w_0_743,w_0_744,w_0_745,w_0_746,w_0_747,w_0_748,w_0_749,w_0_750,w_0_751,w_0_752,w_0_753,w_0_754,w_0_755,w_0_756,w_0_757,w_0_758,w_0_759,w_0_760,w_0_761,w_0_762,w_0_763,w_0_764,w_0_765,w_0_766,w_0_767,w_0_768,w_0_769,w_0_770,w_0_771,w_0_772,w_0_773,w_0_774,w_0_775,w_0_776,w_0_777,w_0_778,w_0_779,w_0_780,w_0_781,w_0_782,w_0_783,w_0_784,
w_1_0,w_1_1,w_1_2,w_1_3,w_1_4,w_1_5,w_1_6,w_1_7,w_1_8,w_1_9,w_1_10,w_1_11,w_1_12,w_1_13,w_1_14,w_1_15,w_1_16,w_1_17,w_1_18,w_1_19,w_1_20,w_1_21,w_1_22,w_1_23,w_1_24,w_1_25,w_1_26,w_1_27,w_1_28,w_1_29,w_1_30,w_1_31,w_1_32,w_1_33,w_1_34,w_1_35,w_1_36,w_1_37,w_1_38,w_1_39,w_1_40,w_1_41,w_1_42,w_1_43,w_1_44,w_1_45,w_1_46,w_1_47,w_1_48,w_1_49,w_1_50,w_1_51,w_1_52,w_1_53,w_1_54,w_1_55,w_1_56,w_1_57,w_1_58,w_1_59,w_1_60,w_1_61,w_1_62,w_1_63,w_1_64,w_1_65,w_1_66,w_1_67,w_1_68,w_1_69,w_1_70,w_1_71,w_1_72,w_1_73,w_1_74,w_1_75,w_1_76,w_1_77,w_1_78,w_1_79,w_1_80,w_1_81,w_1_82,w_1_83,w_1_84,w_1_85,w_1_86,w_1_87,w_1_88,w_1_89,w_1_90,w_1_91,w_1_92,w_1_93,w_1_94,w_1_95,w_1_96,w_1_97,w_1_98,w_1_99,w_1_100,w_1_101,w_1_102,w_1_103,w_1_104,w_1_105,w_1_106,w_1_107,w_1_108,w_1_109,w_1_110,w_1_111,w_1_112,w_1_113,w_1_114,w_1_115,w_1_116,w_1_117,w_1_118,w_1_119,w_1_120,w_1_121,w_1_122,w_1_123,w_1_124,w_1_125,w_1_126,w_1_127,w_1_128,w_1_129,w_1_130,w_1_131,w_1_132,w_1_133,w_1_134,w_1_135,w_1_136,w_1_137,w_1_138,w_1_139,w_1_140,w_1_141,w_1_142,w_1_143,w_1_144,w_1_145,w_1_146,w_1_147,w_1_148,w_1_149,w_1_150,w_1_151,w_1_152,w_1_153,w_1_154,w_1_155,w_1_156,w_1_157,w_1_158,w_1_159,w_1_160,w_1_161,w_1_162,w_1_163,w_1_164,w_1_165,w_1_166,w_1_167,w_1_168,w_1_169,w_1_170,w_1_171,w_1_172,w_1_173,w_1_174,w_1_175,w_1_176,w_1_177,w_1_178,w_1_179,w_1_180,w_1_181,w_1_182,w_1_183,w_1_184,w_1_185,w_1_186,w_1_187,w_1_188,w_1_189,w_1_190,w_1_191,w_1_192,w_1_193,w_1_194,w_1_195,w_1_196,w_1_197,w_1_198,w_1_199,w_1_200,w_1_201,w_1_202,w_1_203,w_1_204,w_1_205,w_1_206,w_1_207,w_1_208,w_1_209,w_1_210,w_1_211,w_1_212,w_1_213,w_1_214,w_1_215,w_1_216,w_1_217,w_1_218,w_1_219,w_1_220,w_1_221,w_1_222,w_1_223,w_1_224,w_1_225,w_1_226,w_1_227,w_1_228,w_1_229,w_1_230,w_1_231,w_1_232,w_1_233,w_1_234,w_1_235,w_1_236,w_1_237,w_1_238,w_1_239,w_1_240,w_1_241,w_1_242,w_1_243,w_1_244,w_1_245,w_1_246,w_1_247,w_1_248,w_1_249,w_1_250,w_1_251,w_1_252,w_1_253,w_1_254,w_1_255,w_1_256,w_1_257,w_1_258,w_1_259,w_1_260,w_1_261,w_1_262,w_1_263,w_1_264,w_1_265,w_1_266,w_1_267,w_1_268,w_1_269,w_1_270,w_1_271,w_1_272,w_1_273,w_1_274,w_1_275,w_1_276,w_1_277,w_1_278,w_1_279,w_1_280,w_1_281,w_1_282,w_1_283,w_1_284,w_1_285,w_1_286,w_1_287,w_1_288,w_1_289,w_1_290,w_1_291,w_1_292,w_1_293,w_1_294,w_1_295,w_1_296,w_1_297,w_1_298,w_1_299,w_1_300,w_1_301,w_1_302,w_1_303,w_1_304,w_1_305,w_1_306,w_1_307,w_1_308,w_1_309,w_1_310,w_1_311,w_1_312,w_1_313,w_1_314,w_1_315,w_1_316,w_1_317,w_1_318,w_1_319,w_1_320,w_1_321,w_1_322,w_1_323,w_1_324,w_1_325,w_1_326,w_1_327,w_1_328,w_1_329,w_1_330,w_1_331,w_1_332,w_1_333,w_1_334,w_1_335,w_1_336,w_1_337,w_1_338,w_1_339,w_1_340,w_1_341,w_1_342,w_1_343,w_1_344,w_1_345,w_1_346,w_1_347,w_1_348,w_1_349,w_1_350,w_1_351,w_1_352,w_1_353,w_1_354,w_1_355,w_1_356,w_1_357,w_1_358,w_1_359,w_1_360,w_1_361,w_1_362,w_1_363,w_1_364,w_1_365,w_1_366,w_1_367,w_1_368,w_1_369,w_1_370,w_1_371,w_1_372,w_1_373,w_1_374,w_1_375,w_1_376,w_1_377,w_1_378,w_1_379,w_1_380,w_1_381,w_1_382,w_1_383,w_1_384,w_1_385,w_1_386,w_1_387,w_1_388,w_1_389,w_1_390,w_1_391,w_1_392,w_1_393,w_1_394,w_1_395,w_1_396,w_1_397,w_1_398,w_1_399,w_1_400,w_1_401,w_1_402,w_1_403,w_1_404,w_1_405,w_1_406,w_1_407,w_1_408,w_1_409,w_1_410,w_1_411,w_1_412,w_1_413,w_1_414,w_1_415,w_1_416,w_1_417,w_1_418,w_1_419,w_1_420,w_1_421,w_1_422,w_1_423,w_1_424,w_1_425,w_1_426,w_1_427,w_1_428,w_1_429,w_1_430,w_1_431,w_1_432,w_1_433,w_1_434,w_1_435,w_1_436,w_1_437,w_1_438,w_1_439,w_1_440,w_1_441,w_1_442,w_1_443,w_1_444,w_1_445,w_1_446,w_1_447,w_1_448,w_1_449,w_1_450,w_1_451,w_1_452,w_1_453,w_1_454,w_1_455,w_1_456,w_1_457,w_1_458,w_1_459,w_1_460,w_1_461,w_1_462,w_1_463,w_1_464,w_1_465,w_1_466,w_1_467,w_1_468,w_1_469,w_1_470,w_1_471,w_1_472,w_1_473,w_1_474,w_1_475,w_1_476,w_1_477,w_1_478,w_1_479,w_1_480,w_1_481,w_1_482,w_1_483,w_1_484,w_1_485,w_1_486,w_1_487,w_1_488,w_1_489,w_1_490,w_1_491,w_1_492,w_1_493,w_1_494,w_1_495,w_1_496,w_1_497,w_1_498,w_1_499,w_1_500,w_1_501,w_1_502,w_1_503,w_1_504,w_1_505,w_1_506,w_1_507,w_1_508,w_1_509,w_1_510,w_1_511,w_1_512,w_1_513,w_1_514,w_1_515,w_1_516,w_1_517,w_1_518,w_1_519,w_1_520,w_1_521,w_1_522,w_1_523,w_1_524,w_1_525,w_1_526,w_1_527,w_1_528,w_1_529,w_1_530,w_1_531,w_1_532,w_1_533,w_1_534,w_1_535,w_1_536,w_1_537,w_1_538,w_1_539,w_1_540,w_1_541,w_1_542,w_1_543,w_1_544,w_1_545,w_1_546,w_1_547,w_1_548,w_1_549,w_1_550,w_1_551,w_1_552,w_1_553,w_1_554,w_1_555,w_1_556,w_1_557,w_1_558,w_1_559,w_1_560,w_1_561,w_1_562,w_1_563,w_1_564,w_1_565,w_1_566,w_1_567,w_1_568,w_1_569,w_1_570,w_1_571,w_1_572,w_1_573,w_1_574,w_1_575,w_1_576,w_1_577,w_1_578,w_1_579,w_1_580,w_1_581,w_1_582,w_1_583,w_1_584,w_1_585,w_1_586,w_1_587,w_1_588,w_1_589,w_1_590,w_1_591,w_1_592,w_1_593,w_1_594,w_1_595,w_1_596,w_1_597,w_1_598,w_1_599,w_1_600,w_1_601,w_1_602,w_1_603,w_1_604,w_1_605,w_1_606,w_1_607,w_1_608,w_1_609,w_1_610,w_1_611,w_1_612,w_1_613,w_1_614,w_1_615,w_1_616,w_1_617,w_1_618,w_1_619,w_1_620,w_1_621,w_1_622,w_1_623,w_1_624,w_1_625,w_1_626,w_1_627,w_1_628,w_1_629,w_1_630,w_1_631,w_1_632,w_1_633,w_1_634,w_1_635,w_1_636,w_1_637,w_1_638,w_1_639,w_1_640,w_1_641,w_1_642,w_1_643,w_1_644,w_1_645,w_1_646,w_1_647,w_1_648,w_1_649,w_1_650,w_1_651,w_1_652,w_1_653,w_1_654,w_1_655,w_1_656,w_1_657,w_1_658,w_1_659,w_1_660,w_1_661,w_1_662,w_1_663,w_1_664,w_1_665,w_1_666,w_1_667,w_1_668,w_1_669,w_1_670,w_1_671,w_1_672,w_1_673,w_1_674,w_1_675,w_1_676,w_1_677,w_1_678,w_1_679,w_1_680,w_1_681,w_1_682,w_1_683,w_1_684,w_1_685,w_1_686,w_1_687,w_1_688,w_1_689,w_1_690,w_1_691,w_1_692,w_1_693,w_1_694,w_1_695,w_1_696,w_1_697,w_1_698,w_1_699,w_1_700,w_1_701,w_1_702,w_1_703,w_1_704,w_1_705,w_1_706,w_1_707,w_1_708,w_1_709,w_1_710,w_1_711,w_1_712,w_1_713,w_1_714,w_1_715,w_1_716,w_1_717,w_1_718,w_1_719,w_1_720,w_1_721,w_1_722,w_1_723,w_1_724,w_1_725,w_1_726,w_1_727,w_1_728,w_1_729,w_1_730,w_1_731,w_1_732,w_1_733,w_1_734,w_1_735,w_1_736,w_1_737,w_1_738,w_1_739,w_1_740,w_1_741,w_1_742,w_1_743,w_1_744,w_1_745,w_1_746,w_1_747,w_1_748,w_1_749,w_1_750,w_1_751,w_1_752,w_1_753,w_1_754,w_1_755,w_1_756,w_1_757,w_1_758,w_1_759,w_1_760,w_1_761,w_1_762,w_1_763,w_1_764,w_1_765,w_1_766,w_1_767,w_1_768,w_1_769,w_1_770,w_1_771,w_1_772,w_1_773,w_1_774,w_1_775,w_1_776,w_1_777,w_1_778,w_1_779,w_1_780,w_1_781,w_1_782,w_1_783,w_1_784,
w_2_0,w_2_1,w_2_2,w_2_3,w_2_4,w_2_5,w_2_6,w_2_7,w_2_8,w_2_9,w_2_10,w_2_11,w_2_12,w_2_13,w_2_14,w_2_15,w_2_16,w_2_17,w_2_18,w_2_19,w_2_20,w_2_21,w_2_22,w_2_23,w_2_24,w_2_25,w_2_26,w_2_27,w_2_28,w_2_29,w_2_30,w_2_31,w_2_32,w_2_33,w_2_34,w_2_35,w_2_36,w_2_37,w_2_38,w_2_39,w_2_40,w_2_41,w_2_42,w_2_43,w_2_44,w_2_45,w_2_46,w_2_47,w_2_48,w_2_49,w_2_50,w_2_51,w_2_52,w_2_53,w_2_54,w_2_55,w_2_56,w_2_57,w_2_58,w_2_59,w_2_60,w_2_61,w_2_62,w_2_63,w_2_64,w_2_65,w_2_66,w_2_67,w_2_68,w_2_69,w_2_70,w_2_71,w_2_72,w_2_73,w_2_74,w_2_75,w_2_76,w_2_77,w_2_78,w_2_79,w_2_80,w_2_81,w_2_82,w_2_83,w_2_84,w_2_85,w_2_86,w_2_87,w_2_88,w_2_89,w_2_90,w_2_91,w_2_92,w_2_93,w_2_94,w_2_95,w_2_96,w_2_97,w_2_98,w_2_99,w_2_100,w_2_101,w_2_102,w_2_103,w_2_104,w_2_105,w_2_106,w_2_107,w_2_108,w_2_109,w_2_110,w_2_111,w_2_112,w_2_113,w_2_114,w_2_115,w_2_116,w_2_117,w_2_118,w_2_119,w_2_120,w_2_121,w_2_122,w_2_123,w_2_124,w_2_125,w_2_126,w_2_127,w_2_128,w_2_129,w_2_130,w_2_131,w_2_132,w_2_133,w_2_134,w_2_135,w_2_136,w_2_137,w_2_138,w_2_139,w_2_140,w_2_141,w_2_142,w_2_143,w_2_144,w_2_145,w_2_146,w_2_147,w_2_148,w_2_149,w_2_150,w_2_151,w_2_152,w_2_153,w_2_154,w_2_155,w_2_156,w_2_157,w_2_158,w_2_159,w_2_160,w_2_161,w_2_162,w_2_163,w_2_164,w_2_165,w_2_166,w_2_167,w_2_168,w_2_169,w_2_170,w_2_171,w_2_172,w_2_173,w_2_174,w_2_175,w_2_176,w_2_177,w_2_178,w_2_179,w_2_180,w_2_181,w_2_182,w_2_183,w_2_184,w_2_185,w_2_186,w_2_187,w_2_188,w_2_189,w_2_190,w_2_191,w_2_192,w_2_193,w_2_194,w_2_195,w_2_196,w_2_197,w_2_198,w_2_199,w_2_200,w_2_201,w_2_202,w_2_203,w_2_204,w_2_205,w_2_206,w_2_207,w_2_208,w_2_209,w_2_210,w_2_211,w_2_212,w_2_213,w_2_214,w_2_215,w_2_216,w_2_217,w_2_218,w_2_219,w_2_220,w_2_221,w_2_222,w_2_223,w_2_224,w_2_225,w_2_226,w_2_227,w_2_228,w_2_229,w_2_230,w_2_231,w_2_232,w_2_233,w_2_234,w_2_235,w_2_236,w_2_237,w_2_238,w_2_239,w_2_240,w_2_241,w_2_242,w_2_243,w_2_244,w_2_245,w_2_246,w_2_247,w_2_248,w_2_249,w_2_250,w_2_251,w_2_252,w_2_253,w_2_254,w_2_255,w_2_256,w_2_257,w_2_258,w_2_259,w_2_260,w_2_261,w_2_262,w_2_263,w_2_264,w_2_265,w_2_266,w_2_267,w_2_268,w_2_269,w_2_270,w_2_271,w_2_272,w_2_273,w_2_274,w_2_275,w_2_276,w_2_277,w_2_278,w_2_279,w_2_280,w_2_281,w_2_282,w_2_283,w_2_284,w_2_285,w_2_286,w_2_287,w_2_288,w_2_289,w_2_290,w_2_291,w_2_292,w_2_293,w_2_294,w_2_295,w_2_296,w_2_297,w_2_298,w_2_299,w_2_300,w_2_301,w_2_302,w_2_303,w_2_304,w_2_305,w_2_306,w_2_307,w_2_308,w_2_309,w_2_310,w_2_311,w_2_312,w_2_313,w_2_314,w_2_315,w_2_316,w_2_317,w_2_318,w_2_319,w_2_320,w_2_321,w_2_322,w_2_323,w_2_324,w_2_325,w_2_326,w_2_327,w_2_328,w_2_329,w_2_330,w_2_331,w_2_332,w_2_333,w_2_334,w_2_335,w_2_336,w_2_337,w_2_338,w_2_339,w_2_340,w_2_341,w_2_342,w_2_343,w_2_344,w_2_345,w_2_346,w_2_347,w_2_348,w_2_349,w_2_350,w_2_351,w_2_352,w_2_353,w_2_354,w_2_355,w_2_356,w_2_357,w_2_358,w_2_359,w_2_360,w_2_361,w_2_362,w_2_363,w_2_364,w_2_365,w_2_366,w_2_367,w_2_368,w_2_369,w_2_370,w_2_371,w_2_372,w_2_373,w_2_374,w_2_375,w_2_376,w_2_377,w_2_378,w_2_379,w_2_380,w_2_381,w_2_382,w_2_383,w_2_384,w_2_385,w_2_386,w_2_387,w_2_388,w_2_389,w_2_390,w_2_391,w_2_392,w_2_393,w_2_394,w_2_395,w_2_396,w_2_397,w_2_398,w_2_399,w_2_400,w_2_401,w_2_402,w_2_403,w_2_404,w_2_405,w_2_406,w_2_407,w_2_408,w_2_409,w_2_410,w_2_411,w_2_412,w_2_413,w_2_414,w_2_415,w_2_416,w_2_417,w_2_418,w_2_419,w_2_420,w_2_421,w_2_422,w_2_423,w_2_424,w_2_425,w_2_426,w_2_427,w_2_428,w_2_429,w_2_430,w_2_431,w_2_432,w_2_433,w_2_434,w_2_435,w_2_436,w_2_437,w_2_438,w_2_439,w_2_440,w_2_441,w_2_442,w_2_443,w_2_444,w_2_445,w_2_446,w_2_447,w_2_448,w_2_449,w_2_450,w_2_451,w_2_452,w_2_453,w_2_454,w_2_455,w_2_456,w_2_457,w_2_458,w_2_459,w_2_460,w_2_461,w_2_462,w_2_463,w_2_464,w_2_465,w_2_466,w_2_467,w_2_468,w_2_469,w_2_470,w_2_471,w_2_472,w_2_473,w_2_474,w_2_475,w_2_476,w_2_477,w_2_478,w_2_479,w_2_480,w_2_481,w_2_482,w_2_483,w_2_484,w_2_485,w_2_486,w_2_487,w_2_488,w_2_489,w_2_490,w_2_491,w_2_492,w_2_493,w_2_494,w_2_495,w_2_496,w_2_497,w_2_498,w_2_499,w_2_500,w_2_501,w_2_502,w_2_503,w_2_504,w_2_505,w_2_506,w_2_507,w_2_508,w_2_509,w_2_510,w_2_511,w_2_512,w_2_513,w_2_514,w_2_515,w_2_516,w_2_517,w_2_518,w_2_519,w_2_520,w_2_521,w_2_522,w_2_523,w_2_524,w_2_525,w_2_526,w_2_527,w_2_528,w_2_529,w_2_530,w_2_531,w_2_532,w_2_533,w_2_534,w_2_535,w_2_536,w_2_537,w_2_538,w_2_539,w_2_540,w_2_541,w_2_542,w_2_543,w_2_544,w_2_545,w_2_546,w_2_547,w_2_548,w_2_549,w_2_550,w_2_551,w_2_552,w_2_553,w_2_554,w_2_555,w_2_556,w_2_557,w_2_558,w_2_559,w_2_560,w_2_561,w_2_562,w_2_563,w_2_564,w_2_565,w_2_566,w_2_567,w_2_568,w_2_569,w_2_570,w_2_571,w_2_572,w_2_573,w_2_574,w_2_575,w_2_576,w_2_577,w_2_578,w_2_579,w_2_580,w_2_581,w_2_582,w_2_583,w_2_584,w_2_585,w_2_586,w_2_587,w_2_588,w_2_589,w_2_590,w_2_591,w_2_592,w_2_593,w_2_594,w_2_595,w_2_596,w_2_597,w_2_598,w_2_599,w_2_600,w_2_601,w_2_602,w_2_603,w_2_604,w_2_605,w_2_606,w_2_607,w_2_608,w_2_609,w_2_610,w_2_611,w_2_612,w_2_613,w_2_614,w_2_615,w_2_616,w_2_617,w_2_618,w_2_619,w_2_620,w_2_621,w_2_622,w_2_623,w_2_624,w_2_625,w_2_626,w_2_627,w_2_628,w_2_629,w_2_630,w_2_631,w_2_632,w_2_633,w_2_634,w_2_635,w_2_636,w_2_637,w_2_638,w_2_639,w_2_640,w_2_641,w_2_642,w_2_643,w_2_644,w_2_645,w_2_646,w_2_647,w_2_648,w_2_649,w_2_650,w_2_651,w_2_652,w_2_653,w_2_654,w_2_655,w_2_656,w_2_657,w_2_658,w_2_659,w_2_660,w_2_661,w_2_662,w_2_663,w_2_664,w_2_665,w_2_666,w_2_667,w_2_668,w_2_669,w_2_670,w_2_671,w_2_672,w_2_673,w_2_674,w_2_675,w_2_676,w_2_677,w_2_678,w_2_679,w_2_680,w_2_681,w_2_682,w_2_683,w_2_684,w_2_685,w_2_686,w_2_687,w_2_688,w_2_689,w_2_690,w_2_691,w_2_692,w_2_693,w_2_694,w_2_695,w_2_696,w_2_697,w_2_698,w_2_699,w_2_700,w_2_701,w_2_702,w_2_703,w_2_704,w_2_705,w_2_706,w_2_707,w_2_708,w_2_709,w_2_710,w_2_711,w_2_712,w_2_713,w_2_714,w_2_715,w_2_716,w_2_717,w_2_718,w_2_719,w_2_720,w_2_721,w_2_722,w_2_723,w_2_724,w_2_725,w_2_726,w_2_727,w_2_728,w_2_729,w_2_730,w_2_731,w_2_732,w_2_733,w_2_734,w_2_735,w_2_736,w_2_737,w_2_738,w_2_739,w_2_740,w_2_741,w_2_742,w_2_743,w_2_744,w_2_745,w_2_746,w_2_747,w_2_748,w_2_749,w_2_750,w_2_751,w_2_752,w_2_753,w_2_754,w_2_755,w_2_756,w_2_757,w_2_758,w_2_759,w_2_760,w_2_761,w_2_762,w_2_763,w_2_764,w_2_765,w_2_766,w_2_767,w_2_768,w_2_769,w_2_770,w_2_771,w_2_772,w_2_773,w_2_774,w_2_775,w_2_776,w_2_777,w_2_778,w_2_779,w_2_780,w_2_781,w_2_782,w_2_783,w_2_784,
w_3_0,w_3_1,w_3_2,w_3_3,w_3_4,w_3_5,w_3_6,w_3_7,w_3_8,w_3_9,w_3_10,w_3_11,w_3_12,w_3_13,w_3_14,w_3_15,w_3_16,w_3_17,w_3_18,w_3_19,w_3_20,w_3_21,w_3_22,w_3_23,w_3_24,w_3_25,w_3_26,w_3_27,w_3_28,w_3_29,w_3_30,w_3_31,w_3_32,w_3_33,w_3_34,w_3_35,w_3_36,w_3_37,w_3_38,w_3_39,w_3_40,w_3_41,w_3_42,w_3_43,w_3_44,w_3_45,w_3_46,w_3_47,w_3_48,w_3_49,w_3_50,w_3_51,w_3_52,w_3_53,w_3_54,w_3_55,w_3_56,w_3_57,w_3_58,w_3_59,w_3_60,w_3_61,w_3_62,w_3_63,w_3_64,w_3_65,w_3_66,w_3_67,w_3_68,w_3_69,w_3_70,w_3_71,w_3_72,w_3_73,w_3_74,w_3_75,w_3_76,w_3_77,w_3_78,w_3_79,w_3_80,w_3_81,w_3_82,w_3_83,w_3_84,w_3_85,w_3_86,w_3_87,w_3_88,w_3_89,w_3_90,w_3_91,w_3_92,w_3_93,w_3_94,w_3_95,w_3_96,w_3_97,w_3_98,w_3_99,w_3_100,w_3_101,w_3_102,w_3_103,w_3_104,w_3_105,w_3_106,w_3_107,w_3_108,w_3_109,w_3_110,w_3_111,w_3_112,w_3_113,w_3_114,w_3_115,w_3_116,w_3_117,w_3_118,w_3_119,w_3_120,w_3_121,w_3_122,w_3_123,w_3_124,w_3_125,w_3_126,w_3_127,w_3_128,w_3_129,w_3_130,w_3_131,w_3_132,w_3_133,w_3_134,w_3_135,w_3_136,w_3_137,w_3_138,w_3_139,w_3_140,w_3_141,w_3_142,w_3_143,w_3_144,w_3_145,w_3_146,w_3_147,w_3_148,w_3_149,w_3_150,w_3_151,w_3_152,w_3_153,w_3_154,w_3_155,w_3_156,w_3_157,w_3_158,w_3_159,w_3_160,w_3_161,w_3_162,w_3_163,w_3_164,w_3_165,w_3_166,w_3_167,w_3_168,w_3_169,w_3_170,w_3_171,w_3_172,w_3_173,w_3_174,w_3_175,w_3_176,w_3_177,w_3_178,w_3_179,w_3_180,w_3_181,w_3_182,w_3_183,w_3_184,w_3_185,w_3_186,w_3_187,w_3_188,w_3_189,w_3_190,w_3_191,w_3_192,w_3_193,w_3_194,w_3_195,w_3_196,w_3_197,w_3_198,w_3_199,w_3_200,w_3_201,w_3_202,w_3_203,w_3_204,w_3_205,w_3_206,w_3_207,w_3_208,w_3_209,w_3_210,w_3_211,w_3_212,w_3_213,w_3_214,w_3_215,w_3_216,w_3_217,w_3_218,w_3_219,w_3_220,w_3_221,w_3_222,w_3_223,w_3_224,w_3_225,w_3_226,w_3_227,w_3_228,w_3_229,w_3_230,w_3_231,w_3_232,w_3_233,w_3_234,w_3_235,w_3_236,w_3_237,w_3_238,w_3_239,w_3_240,w_3_241,w_3_242,w_3_243,w_3_244,w_3_245,w_3_246,w_3_247,w_3_248,w_3_249,w_3_250,w_3_251,w_3_252,w_3_253,w_3_254,w_3_255,w_3_256,w_3_257,w_3_258,w_3_259,w_3_260,w_3_261,w_3_262,w_3_263,w_3_264,w_3_265,w_3_266,w_3_267,w_3_268,w_3_269,w_3_270,w_3_271,w_3_272,w_3_273,w_3_274,w_3_275,w_3_276,w_3_277,w_3_278,w_3_279,w_3_280,w_3_281,w_3_282,w_3_283,w_3_284,w_3_285,w_3_286,w_3_287,w_3_288,w_3_289,w_3_290,w_3_291,w_3_292,w_3_293,w_3_294,w_3_295,w_3_296,w_3_297,w_3_298,w_3_299,w_3_300,w_3_301,w_3_302,w_3_303,w_3_304,w_3_305,w_3_306,w_3_307,w_3_308,w_3_309,w_3_310,w_3_311,w_3_312,w_3_313,w_3_314,w_3_315,w_3_316,w_3_317,w_3_318,w_3_319,w_3_320,w_3_321,w_3_322,w_3_323,w_3_324,w_3_325,w_3_326,w_3_327,w_3_328,w_3_329,w_3_330,w_3_331,w_3_332,w_3_333,w_3_334,w_3_335,w_3_336,w_3_337,w_3_338,w_3_339,w_3_340,w_3_341,w_3_342,w_3_343,w_3_344,w_3_345,w_3_346,w_3_347,w_3_348,w_3_349,w_3_350,w_3_351,w_3_352,w_3_353,w_3_354,w_3_355,w_3_356,w_3_357,w_3_358,w_3_359,w_3_360,w_3_361,w_3_362,w_3_363,w_3_364,w_3_365,w_3_366,w_3_367,w_3_368,w_3_369,w_3_370,w_3_371,w_3_372,w_3_373,w_3_374,w_3_375,w_3_376,w_3_377,w_3_378,w_3_379,w_3_380,w_3_381,w_3_382,w_3_383,w_3_384,w_3_385,w_3_386,w_3_387,w_3_388,w_3_389,w_3_390,w_3_391,w_3_392,w_3_393,w_3_394,w_3_395,w_3_396,w_3_397,w_3_398,w_3_399,w_3_400,w_3_401,w_3_402,w_3_403,w_3_404,w_3_405,w_3_406,w_3_407,w_3_408,w_3_409,w_3_410,w_3_411,w_3_412,w_3_413,w_3_414,w_3_415,w_3_416,w_3_417,w_3_418,w_3_419,w_3_420,w_3_421,w_3_422,w_3_423,w_3_424,w_3_425,w_3_426,w_3_427,w_3_428,w_3_429,w_3_430,w_3_431,w_3_432,w_3_433,w_3_434,w_3_435,w_3_436,w_3_437,w_3_438,w_3_439,w_3_440,w_3_441,w_3_442,w_3_443,w_3_444,w_3_445,w_3_446,w_3_447,w_3_448,w_3_449,w_3_450,w_3_451,w_3_452,w_3_453,w_3_454,w_3_455,w_3_456,w_3_457,w_3_458,w_3_459,w_3_460,w_3_461,w_3_462,w_3_463,w_3_464,w_3_465,w_3_466,w_3_467,w_3_468,w_3_469,w_3_470,w_3_471,w_3_472,w_3_473,w_3_474,w_3_475,w_3_476,w_3_477,w_3_478,w_3_479,w_3_480,w_3_481,w_3_482,w_3_483,w_3_484,w_3_485,w_3_486,w_3_487,w_3_488,w_3_489,w_3_490,w_3_491,w_3_492,w_3_493,w_3_494,w_3_495,w_3_496,w_3_497,w_3_498,w_3_499,w_3_500,w_3_501,w_3_502,w_3_503,w_3_504,w_3_505,w_3_506,w_3_507,w_3_508,w_3_509,w_3_510,w_3_511,w_3_512,w_3_513,w_3_514,w_3_515,w_3_516,w_3_517,w_3_518,w_3_519,w_3_520,w_3_521,w_3_522,w_3_523,w_3_524,w_3_525,w_3_526,w_3_527,w_3_528,w_3_529,w_3_530,w_3_531,w_3_532,w_3_533,w_3_534,w_3_535,w_3_536,w_3_537,w_3_538,w_3_539,w_3_540,w_3_541,w_3_542,w_3_543,w_3_544,w_3_545,w_3_546,w_3_547,w_3_548,w_3_549,w_3_550,w_3_551,w_3_552,w_3_553,w_3_554,w_3_555,w_3_556,w_3_557,w_3_558,w_3_559,w_3_560,w_3_561,w_3_562,w_3_563,w_3_564,w_3_565,w_3_566,w_3_567,w_3_568,w_3_569,w_3_570,w_3_571,w_3_572,w_3_573,w_3_574,w_3_575,w_3_576,w_3_577,w_3_578,w_3_579,w_3_580,w_3_581,w_3_582,w_3_583,w_3_584,w_3_585,w_3_586,w_3_587,w_3_588,w_3_589,w_3_590,w_3_591,w_3_592,w_3_593,w_3_594,w_3_595,w_3_596,w_3_597,w_3_598,w_3_599,w_3_600,w_3_601,w_3_602,w_3_603,w_3_604,w_3_605,w_3_606,w_3_607,w_3_608,w_3_609,w_3_610,w_3_611,w_3_612,w_3_613,w_3_614,w_3_615,w_3_616,w_3_617,w_3_618,w_3_619,w_3_620,w_3_621,w_3_622,w_3_623,w_3_624,w_3_625,w_3_626,w_3_627,w_3_628,w_3_629,w_3_630,w_3_631,w_3_632,w_3_633,w_3_634,w_3_635,w_3_636,w_3_637,w_3_638,w_3_639,w_3_640,w_3_641,w_3_642,w_3_643,w_3_644,w_3_645,w_3_646,w_3_647,w_3_648,w_3_649,w_3_650,w_3_651,w_3_652,w_3_653,w_3_654,w_3_655,w_3_656,w_3_657,w_3_658,w_3_659,w_3_660,w_3_661,w_3_662,w_3_663,w_3_664,w_3_665,w_3_666,w_3_667,w_3_668,w_3_669,w_3_670,w_3_671,w_3_672,w_3_673,w_3_674,w_3_675,w_3_676,w_3_677,w_3_678,w_3_679,w_3_680,w_3_681,w_3_682,w_3_683,w_3_684,w_3_685,w_3_686,w_3_687,w_3_688,w_3_689,w_3_690,w_3_691,w_3_692,w_3_693,w_3_694,w_3_695,w_3_696,w_3_697,w_3_698,w_3_699,w_3_700,w_3_701,w_3_702,w_3_703,w_3_704,w_3_705,w_3_706,w_3_707,w_3_708,w_3_709,w_3_710,w_3_711,w_3_712,w_3_713,w_3_714,w_3_715,w_3_716,w_3_717,w_3_718,w_3_719,w_3_720,w_3_721,w_3_722,w_3_723,w_3_724,w_3_725,w_3_726,w_3_727,w_3_728,w_3_729,w_3_730,w_3_731,w_3_732,w_3_733,w_3_734,w_3_735,w_3_736,w_3_737,w_3_738,w_3_739,w_3_740,w_3_741,w_3_742,w_3_743,w_3_744,w_3_745,w_3_746,w_3_747,w_3_748,w_3_749,w_3_750,w_3_751,w_3_752,w_3_753,w_3_754,w_3_755,w_3_756,w_3_757,w_3_758,w_3_759,w_3_760,w_3_761,w_3_762,w_3_763,w_3_764,w_3_765,w_3_766,w_3_767,w_3_768,w_3_769,w_3_770,w_3_771,w_3_772,w_3_773,w_3_774,w_3_775,w_3_776,w_3_777,w_3_778,w_3_779,w_3_780,w_3_781,w_3_782,w_3_783,w_3_784,
w_4_0,w_4_1,w_4_2,w_4_3,w_4_4,w_4_5,w_4_6,w_4_7,w_4_8,w_4_9,w_4_10,w_4_11,w_4_12,w_4_13,w_4_14,w_4_15,w_4_16,w_4_17,w_4_18,w_4_19,w_4_20,w_4_21,w_4_22,w_4_23,w_4_24,w_4_25,w_4_26,w_4_27,w_4_28,w_4_29,w_4_30,w_4_31,w_4_32,w_4_33,w_4_34,w_4_35,w_4_36,w_4_37,w_4_38,w_4_39,w_4_40,w_4_41,w_4_42,w_4_43,w_4_44,w_4_45,w_4_46,w_4_47,w_4_48,w_4_49,w_4_50,w_4_51,w_4_52,w_4_53,w_4_54,w_4_55,w_4_56,w_4_57,w_4_58,w_4_59,w_4_60,w_4_61,w_4_62,w_4_63,w_4_64,w_4_65,w_4_66,w_4_67,w_4_68,w_4_69,w_4_70,w_4_71,w_4_72,w_4_73,w_4_74,w_4_75,w_4_76,w_4_77,w_4_78,w_4_79,w_4_80,w_4_81,w_4_82,w_4_83,w_4_84,w_4_85,w_4_86,w_4_87,w_4_88,w_4_89,w_4_90,w_4_91,w_4_92,w_4_93,w_4_94,w_4_95,w_4_96,w_4_97,w_4_98,w_4_99,w_4_100,w_4_101,w_4_102,w_4_103,w_4_104,w_4_105,w_4_106,w_4_107,w_4_108,w_4_109,w_4_110,w_4_111,w_4_112,w_4_113,w_4_114,w_4_115,w_4_116,w_4_117,w_4_118,w_4_119,w_4_120,w_4_121,w_4_122,w_4_123,w_4_124,w_4_125,w_4_126,w_4_127,w_4_128,w_4_129,w_4_130,w_4_131,w_4_132,w_4_133,w_4_134,w_4_135,w_4_136,w_4_137,w_4_138,w_4_139,w_4_140,w_4_141,w_4_142,w_4_143,w_4_144,w_4_145,w_4_146,w_4_147,w_4_148,w_4_149,w_4_150,w_4_151,w_4_152,w_4_153,w_4_154,w_4_155,w_4_156,w_4_157,w_4_158,w_4_159,w_4_160,w_4_161,w_4_162,w_4_163,w_4_164,w_4_165,w_4_166,w_4_167,w_4_168,w_4_169,w_4_170,w_4_171,w_4_172,w_4_173,w_4_174,w_4_175,w_4_176,w_4_177,w_4_178,w_4_179,w_4_180,w_4_181,w_4_182,w_4_183,w_4_184,w_4_185,w_4_186,w_4_187,w_4_188,w_4_189,w_4_190,w_4_191,w_4_192,w_4_193,w_4_194,w_4_195,w_4_196,w_4_197,w_4_198,w_4_199,w_4_200,w_4_201,w_4_202,w_4_203,w_4_204,w_4_205,w_4_206,w_4_207,w_4_208,w_4_209,w_4_210,w_4_211,w_4_212,w_4_213,w_4_214,w_4_215,w_4_216,w_4_217,w_4_218,w_4_219,w_4_220,w_4_221,w_4_222,w_4_223,w_4_224,w_4_225,w_4_226,w_4_227,w_4_228,w_4_229,w_4_230,w_4_231,w_4_232,w_4_233,w_4_234,w_4_235,w_4_236,w_4_237,w_4_238,w_4_239,w_4_240,w_4_241,w_4_242,w_4_243,w_4_244,w_4_245,w_4_246,w_4_247,w_4_248,w_4_249,w_4_250,w_4_251,w_4_252,w_4_253,w_4_254,w_4_255,w_4_256,w_4_257,w_4_258,w_4_259,w_4_260,w_4_261,w_4_262,w_4_263,w_4_264,w_4_265,w_4_266,w_4_267,w_4_268,w_4_269,w_4_270,w_4_271,w_4_272,w_4_273,w_4_274,w_4_275,w_4_276,w_4_277,w_4_278,w_4_279,w_4_280,w_4_281,w_4_282,w_4_283,w_4_284,w_4_285,w_4_286,w_4_287,w_4_288,w_4_289,w_4_290,w_4_291,w_4_292,w_4_293,w_4_294,w_4_295,w_4_296,w_4_297,w_4_298,w_4_299,w_4_300,w_4_301,w_4_302,w_4_303,w_4_304,w_4_305,w_4_306,w_4_307,w_4_308,w_4_309,w_4_310,w_4_311,w_4_312,w_4_313,w_4_314,w_4_315,w_4_316,w_4_317,w_4_318,w_4_319,w_4_320,w_4_321,w_4_322,w_4_323,w_4_324,w_4_325,w_4_326,w_4_327,w_4_328,w_4_329,w_4_330,w_4_331,w_4_332,w_4_333,w_4_334,w_4_335,w_4_336,w_4_337,w_4_338,w_4_339,w_4_340,w_4_341,w_4_342,w_4_343,w_4_344,w_4_345,w_4_346,w_4_347,w_4_348,w_4_349,w_4_350,w_4_351,w_4_352,w_4_353,w_4_354,w_4_355,w_4_356,w_4_357,w_4_358,w_4_359,w_4_360,w_4_361,w_4_362,w_4_363,w_4_364,w_4_365,w_4_366,w_4_367,w_4_368,w_4_369,w_4_370,w_4_371,w_4_372,w_4_373,w_4_374,w_4_375,w_4_376,w_4_377,w_4_378,w_4_379,w_4_380,w_4_381,w_4_382,w_4_383,w_4_384,w_4_385,w_4_386,w_4_387,w_4_388,w_4_389,w_4_390,w_4_391,w_4_392,w_4_393,w_4_394,w_4_395,w_4_396,w_4_397,w_4_398,w_4_399,w_4_400,w_4_401,w_4_402,w_4_403,w_4_404,w_4_405,w_4_406,w_4_407,w_4_408,w_4_409,w_4_410,w_4_411,w_4_412,w_4_413,w_4_414,w_4_415,w_4_416,w_4_417,w_4_418,w_4_419,w_4_420,w_4_421,w_4_422,w_4_423,w_4_424,w_4_425,w_4_426,w_4_427,w_4_428,w_4_429,w_4_430,w_4_431,w_4_432,w_4_433,w_4_434,w_4_435,w_4_436,w_4_437,w_4_438,w_4_439,w_4_440,w_4_441,w_4_442,w_4_443,w_4_444,w_4_445,w_4_446,w_4_447,w_4_448,w_4_449,w_4_450,w_4_451,w_4_452,w_4_453,w_4_454,w_4_455,w_4_456,w_4_457,w_4_458,w_4_459,w_4_460,w_4_461,w_4_462,w_4_463,w_4_464,w_4_465,w_4_466,w_4_467,w_4_468,w_4_469,w_4_470,w_4_471,w_4_472,w_4_473,w_4_474,w_4_475,w_4_476,w_4_477,w_4_478,w_4_479,w_4_480,w_4_481,w_4_482,w_4_483,w_4_484,w_4_485,w_4_486,w_4_487,w_4_488,w_4_489,w_4_490,w_4_491,w_4_492,w_4_493,w_4_494,w_4_495,w_4_496,w_4_497,w_4_498,w_4_499,w_4_500,w_4_501,w_4_502,w_4_503,w_4_504,w_4_505,w_4_506,w_4_507,w_4_508,w_4_509,w_4_510,w_4_511,w_4_512,w_4_513,w_4_514,w_4_515,w_4_516,w_4_517,w_4_518,w_4_519,w_4_520,w_4_521,w_4_522,w_4_523,w_4_524,w_4_525,w_4_526,w_4_527,w_4_528,w_4_529,w_4_530,w_4_531,w_4_532,w_4_533,w_4_534,w_4_535,w_4_536,w_4_537,w_4_538,w_4_539,w_4_540,w_4_541,w_4_542,w_4_543,w_4_544,w_4_545,w_4_546,w_4_547,w_4_548,w_4_549,w_4_550,w_4_551,w_4_552,w_4_553,w_4_554,w_4_555,w_4_556,w_4_557,w_4_558,w_4_559,w_4_560,w_4_561,w_4_562,w_4_563,w_4_564,w_4_565,w_4_566,w_4_567,w_4_568,w_4_569,w_4_570,w_4_571,w_4_572,w_4_573,w_4_574,w_4_575,w_4_576,w_4_577,w_4_578,w_4_579,w_4_580,w_4_581,w_4_582,w_4_583,w_4_584,w_4_585,w_4_586,w_4_587,w_4_588,w_4_589,w_4_590,w_4_591,w_4_592,w_4_593,w_4_594,w_4_595,w_4_596,w_4_597,w_4_598,w_4_599,w_4_600,w_4_601,w_4_602,w_4_603,w_4_604,w_4_605,w_4_606,w_4_607,w_4_608,w_4_609,w_4_610,w_4_611,w_4_612,w_4_613,w_4_614,w_4_615,w_4_616,w_4_617,w_4_618,w_4_619,w_4_620,w_4_621,w_4_622,w_4_623,w_4_624,w_4_625,w_4_626,w_4_627,w_4_628,w_4_629,w_4_630,w_4_631,w_4_632,w_4_633,w_4_634,w_4_635,w_4_636,w_4_637,w_4_638,w_4_639,w_4_640,w_4_641,w_4_642,w_4_643,w_4_644,w_4_645,w_4_646,w_4_647,w_4_648,w_4_649,w_4_650,w_4_651,w_4_652,w_4_653,w_4_654,w_4_655,w_4_656,w_4_657,w_4_658,w_4_659,w_4_660,w_4_661,w_4_662,w_4_663,w_4_664,w_4_665,w_4_666,w_4_667,w_4_668,w_4_669,w_4_670,w_4_671,w_4_672,w_4_673,w_4_674,w_4_675,w_4_676,w_4_677,w_4_678,w_4_679,w_4_680,w_4_681,w_4_682,w_4_683,w_4_684,w_4_685,w_4_686,w_4_687,w_4_688,w_4_689,w_4_690,w_4_691,w_4_692,w_4_693,w_4_694,w_4_695,w_4_696,w_4_697,w_4_698,w_4_699,w_4_700,w_4_701,w_4_702,w_4_703,w_4_704,w_4_705,w_4_706,w_4_707,w_4_708,w_4_709,w_4_710,w_4_711,w_4_712,w_4_713,w_4_714,w_4_715,w_4_716,w_4_717,w_4_718,w_4_719,w_4_720,w_4_721,w_4_722,w_4_723,w_4_724,w_4_725,w_4_726,w_4_727,w_4_728,w_4_729,w_4_730,w_4_731,w_4_732,w_4_733,w_4_734,w_4_735,w_4_736,w_4_737,w_4_738,w_4_739,w_4_740,w_4_741,w_4_742,w_4_743,w_4_744,w_4_745,w_4_746,w_4_747,w_4_748,w_4_749,w_4_750,w_4_751,w_4_752,w_4_753,w_4_754,w_4_755,w_4_756,w_4_757,w_4_758,w_4_759,w_4_760,w_4_761,w_4_762,w_4_763,w_4_764,w_4_765,w_4_766,w_4_767,w_4_768,w_4_769,w_4_770,w_4_771,w_4_772,w_4_773,w_4_774,w_4_775,w_4_776,w_4_777,w_4_778,w_4_779,w_4_780,w_4_781,w_4_782,w_4_783,w_4_784,
w_5_0,w_5_1,w_5_2,w_5_3,w_5_4,w_5_5,w_5_6,w_5_7,w_5_8,w_5_9,w_5_10,w_5_11,w_5_12,w_5_13,w_5_14,w_5_15,w_5_16,w_5_17,w_5_18,w_5_19,w_5_20,w_5_21,w_5_22,w_5_23,w_5_24,w_5_25,w_5_26,w_5_27,w_5_28,w_5_29,w_5_30,w_5_31,w_5_32,w_5_33,w_5_34,w_5_35,w_5_36,w_5_37,w_5_38,w_5_39,w_5_40,w_5_41,w_5_42,w_5_43,w_5_44,w_5_45,w_5_46,w_5_47,w_5_48,w_5_49,w_5_50,w_5_51,w_5_52,w_5_53,w_5_54,w_5_55,w_5_56,w_5_57,w_5_58,w_5_59,w_5_60,w_5_61,w_5_62,w_5_63,w_5_64,w_5_65,w_5_66,w_5_67,w_5_68,w_5_69,w_5_70,w_5_71,w_5_72,w_5_73,w_5_74,w_5_75,w_5_76,w_5_77,w_5_78,w_5_79,w_5_80,w_5_81,w_5_82,w_5_83,w_5_84,w_5_85,w_5_86,w_5_87,w_5_88,w_5_89,w_5_90,w_5_91,w_5_92,w_5_93,w_5_94,w_5_95,w_5_96,w_5_97,w_5_98,w_5_99,w_5_100,w_5_101,w_5_102,w_5_103,w_5_104,w_5_105,w_5_106,w_5_107,w_5_108,w_5_109,w_5_110,w_5_111,w_5_112,w_5_113,w_5_114,w_5_115,w_5_116,w_5_117,w_5_118,w_5_119,w_5_120,w_5_121,w_5_122,w_5_123,w_5_124,w_5_125,w_5_126,w_5_127,w_5_128,w_5_129,w_5_130,w_5_131,w_5_132,w_5_133,w_5_134,w_5_135,w_5_136,w_5_137,w_5_138,w_5_139,w_5_140,w_5_141,w_5_142,w_5_143,w_5_144,w_5_145,w_5_146,w_5_147,w_5_148,w_5_149,w_5_150,w_5_151,w_5_152,w_5_153,w_5_154,w_5_155,w_5_156,w_5_157,w_5_158,w_5_159,w_5_160,w_5_161,w_5_162,w_5_163,w_5_164,w_5_165,w_5_166,w_5_167,w_5_168,w_5_169,w_5_170,w_5_171,w_5_172,w_5_173,w_5_174,w_5_175,w_5_176,w_5_177,w_5_178,w_5_179,w_5_180,w_5_181,w_5_182,w_5_183,w_5_184,w_5_185,w_5_186,w_5_187,w_5_188,w_5_189,w_5_190,w_5_191,w_5_192,w_5_193,w_5_194,w_5_195,w_5_196,w_5_197,w_5_198,w_5_199,w_5_200,w_5_201,w_5_202,w_5_203,w_5_204,w_5_205,w_5_206,w_5_207,w_5_208,w_5_209,w_5_210,w_5_211,w_5_212,w_5_213,w_5_214,w_5_215,w_5_216,w_5_217,w_5_218,w_5_219,w_5_220,w_5_221,w_5_222,w_5_223,w_5_224,w_5_225,w_5_226,w_5_227,w_5_228,w_5_229,w_5_230,w_5_231,w_5_232,w_5_233,w_5_234,w_5_235,w_5_236,w_5_237,w_5_238,w_5_239,w_5_240,w_5_241,w_5_242,w_5_243,w_5_244,w_5_245,w_5_246,w_5_247,w_5_248,w_5_249,w_5_250,w_5_251,w_5_252,w_5_253,w_5_254,w_5_255,w_5_256,w_5_257,w_5_258,w_5_259,w_5_260,w_5_261,w_5_262,w_5_263,w_5_264,w_5_265,w_5_266,w_5_267,w_5_268,w_5_269,w_5_270,w_5_271,w_5_272,w_5_273,w_5_274,w_5_275,w_5_276,w_5_277,w_5_278,w_5_279,w_5_280,w_5_281,w_5_282,w_5_283,w_5_284,w_5_285,w_5_286,w_5_287,w_5_288,w_5_289,w_5_290,w_5_291,w_5_292,w_5_293,w_5_294,w_5_295,w_5_296,w_5_297,w_5_298,w_5_299,w_5_300,w_5_301,w_5_302,w_5_303,w_5_304,w_5_305,w_5_306,w_5_307,w_5_308,w_5_309,w_5_310,w_5_311,w_5_312,w_5_313,w_5_314,w_5_315,w_5_316,w_5_317,w_5_318,w_5_319,w_5_320,w_5_321,w_5_322,w_5_323,w_5_324,w_5_325,w_5_326,w_5_327,w_5_328,w_5_329,w_5_330,w_5_331,w_5_332,w_5_333,w_5_334,w_5_335,w_5_336,w_5_337,w_5_338,w_5_339,w_5_340,w_5_341,w_5_342,w_5_343,w_5_344,w_5_345,w_5_346,w_5_347,w_5_348,w_5_349,w_5_350,w_5_351,w_5_352,w_5_353,w_5_354,w_5_355,w_5_356,w_5_357,w_5_358,w_5_359,w_5_360,w_5_361,w_5_362,w_5_363,w_5_364,w_5_365,w_5_366,w_5_367,w_5_368,w_5_369,w_5_370,w_5_371,w_5_372,w_5_373,w_5_374,w_5_375,w_5_376,w_5_377,w_5_378,w_5_379,w_5_380,w_5_381,w_5_382,w_5_383,w_5_384,w_5_385,w_5_386,w_5_387,w_5_388,w_5_389,w_5_390,w_5_391,w_5_392,w_5_393,w_5_394,w_5_395,w_5_396,w_5_397,w_5_398,w_5_399,w_5_400,w_5_401,w_5_402,w_5_403,w_5_404,w_5_405,w_5_406,w_5_407,w_5_408,w_5_409,w_5_410,w_5_411,w_5_412,w_5_413,w_5_414,w_5_415,w_5_416,w_5_417,w_5_418,w_5_419,w_5_420,w_5_421,w_5_422,w_5_423,w_5_424,w_5_425,w_5_426,w_5_427,w_5_428,w_5_429,w_5_430,w_5_431,w_5_432,w_5_433,w_5_434,w_5_435,w_5_436,w_5_437,w_5_438,w_5_439,w_5_440,w_5_441,w_5_442,w_5_443,w_5_444,w_5_445,w_5_446,w_5_447,w_5_448,w_5_449,w_5_450,w_5_451,w_5_452,w_5_453,w_5_454,w_5_455,w_5_456,w_5_457,w_5_458,w_5_459,w_5_460,w_5_461,w_5_462,w_5_463,w_5_464,w_5_465,w_5_466,w_5_467,w_5_468,w_5_469,w_5_470,w_5_471,w_5_472,w_5_473,w_5_474,w_5_475,w_5_476,w_5_477,w_5_478,w_5_479,w_5_480,w_5_481,w_5_482,w_5_483,w_5_484,w_5_485,w_5_486,w_5_487,w_5_488,w_5_489,w_5_490,w_5_491,w_5_492,w_5_493,w_5_494,w_5_495,w_5_496,w_5_497,w_5_498,w_5_499,w_5_500,w_5_501,w_5_502,w_5_503,w_5_504,w_5_505,w_5_506,w_5_507,w_5_508,w_5_509,w_5_510,w_5_511,w_5_512,w_5_513,w_5_514,w_5_515,w_5_516,w_5_517,w_5_518,w_5_519,w_5_520,w_5_521,w_5_522,w_5_523,w_5_524,w_5_525,w_5_526,w_5_527,w_5_528,w_5_529,w_5_530,w_5_531,w_5_532,w_5_533,w_5_534,w_5_535,w_5_536,w_5_537,w_5_538,w_5_539,w_5_540,w_5_541,w_5_542,w_5_543,w_5_544,w_5_545,w_5_546,w_5_547,w_5_548,w_5_549,w_5_550,w_5_551,w_5_552,w_5_553,w_5_554,w_5_555,w_5_556,w_5_557,w_5_558,w_5_559,w_5_560,w_5_561,w_5_562,w_5_563,w_5_564,w_5_565,w_5_566,w_5_567,w_5_568,w_5_569,w_5_570,w_5_571,w_5_572,w_5_573,w_5_574,w_5_575,w_5_576,w_5_577,w_5_578,w_5_579,w_5_580,w_5_581,w_5_582,w_5_583,w_5_584,w_5_585,w_5_586,w_5_587,w_5_588,w_5_589,w_5_590,w_5_591,w_5_592,w_5_593,w_5_594,w_5_595,w_5_596,w_5_597,w_5_598,w_5_599,w_5_600,w_5_601,w_5_602,w_5_603,w_5_604,w_5_605,w_5_606,w_5_607,w_5_608,w_5_609,w_5_610,w_5_611,w_5_612,w_5_613,w_5_614,w_5_615,w_5_616,w_5_617,w_5_618,w_5_619,w_5_620,w_5_621,w_5_622,w_5_623,w_5_624,w_5_625,w_5_626,w_5_627,w_5_628,w_5_629,w_5_630,w_5_631,w_5_632,w_5_633,w_5_634,w_5_635,w_5_636,w_5_637,w_5_638,w_5_639,w_5_640,w_5_641,w_5_642,w_5_643,w_5_644,w_5_645,w_5_646,w_5_647,w_5_648,w_5_649,w_5_650,w_5_651,w_5_652,w_5_653,w_5_654,w_5_655,w_5_656,w_5_657,w_5_658,w_5_659,w_5_660,w_5_661,w_5_662,w_5_663,w_5_664,w_5_665,w_5_666,w_5_667,w_5_668,w_5_669,w_5_670,w_5_671,w_5_672,w_5_673,w_5_674,w_5_675,w_5_676,w_5_677,w_5_678,w_5_679,w_5_680,w_5_681,w_5_682,w_5_683,w_5_684,w_5_685,w_5_686,w_5_687,w_5_688,w_5_689,w_5_690,w_5_691,w_5_692,w_5_693,w_5_694,w_5_695,w_5_696,w_5_697,w_5_698,w_5_699,w_5_700,w_5_701,w_5_702,w_5_703,w_5_704,w_5_705,w_5_706,w_5_707,w_5_708,w_5_709,w_5_710,w_5_711,w_5_712,w_5_713,w_5_714,w_5_715,w_5_716,w_5_717,w_5_718,w_5_719,w_5_720,w_5_721,w_5_722,w_5_723,w_5_724,w_5_725,w_5_726,w_5_727,w_5_728,w_5_729,w_5_730,w_5_731,w_5_732,w_5_733,w_5_734,w_5_735,w_5_736,w_5_737,w_5_738,w_5_739,w_5_740,w_5_741,w_5_742,w_5_743,w_5_744,w_5_745,w_5_746,w_5_747,w_5_748,w_5_749,w_5_750,w_5_751,w_5_752,w_5_753,w_5_754,w_5_755,w_5_756,w_5_757,w_5_758,w_5_759,w_5_760,w_5_761,w_5_762,w_5_763,w_5_764,w_5_765,w_5_766,w_5_767,w_5_768,w_5_769,w_5_770,w_5_771,w_5_772,w_5_773,w_5_774,w_5_775,w_5_776,w_5_777,w_5_778,w_5_779,w_5_780,w_5_781,w_5_782,w_5_783,w_5_784,
w_6_0,w_6_1,w_6_2,w_6_3,w_6_4,w_6_5,w_6_6,w_6_7,w_6_8,w_6_9,w_6_10,w_6_11,w_6_12,w_6_13,w_6_14,w_6_15,w_6_16,w_6_17,w_6_18,w_6_19,w_6_20,w_6_21,w_6_22,w_6_23,w_6_24,w_6_25,w_6_26,w_6_27,w_6_28,w_6_29,w_6_30,w_6_31,w_6_32,w_6_33,w_6_34,w_6_35,w_6_36,w_6_37,w_6_38,w_6_39,w_6_40,w_6_41,w_6_42,w_6_43,w_6_44,w_6_45,w_6_46,w_6_47,w_6_48,w_6_49,w_6_50,w_6_51,w_6_52,w_6_53,w_6_54,w_6_55,w_6_56,w_6_57,w_6_58,w_6_59,w_6_60,w_6_61,w_6_62,w_6_63,w_6_64,w_6_65,w_6_66,w_6_67,w_6_68,w_6_69,w_6_70,w_6_71,w_6_72,w_6_73,w_6_74,w_6_75,w_6_76,w_6_77,w_6_78,w_6_79,w_6_80,w_6_81,w_6_82,w_6_83,w_6_84,w_6_85,w_6_86,w_6_87,w_6_88,w_6_89,w_6_90,w_6_91,w_6_92,w_6_93,w_6_94,w_6_95,w_6_96,w_6_97,w_6_98,w_6_99,w_6_100,w_6_101,w_6_102,w_6_103,w_6_104,w_6_105,w_6_106,w_6_107,w_6_108,w_6_109,w_6_110,w_6_111,w_6_112,w_6_113,w_6_114,w_6_115,w_6_116,w_6_117,w_6_118,w_6_119,w_6_120,w_6_121,w_6_122,w_6_123,w_6_124,w_6_125,w_6_126,w_6_127,w_6_128,w_6_129,w_6_130,w_6_131,w_6_132,w_6_133,w_6_134,w_6_135,w_6_136,w_6_137,w_6_138,w_6_139,w_6_140,w_6_141,w_6_142,w_6_143,w_6_144,w_6_145,w_6_146,w_6_147,w_6_148,w_6_149,w_6_150,w_6_151,w_6_152,w_6_153,w_6_154,w_6_155,w_6_156,w_6_157,w_6_158,w_6_159,w_6_160,w_6_161,w_6_162,w_6_163,w_6_164,w_6_165,w_6_166,w_6_167,w_6_168,w_6_169,w_6_170,w_6_171,w_6_172,w_6_173,w_6_174,w_6_175,w_6_176,w_6_177,w_6_178,w_6_179,w_6_180,w_6_181,w_6_182,w_6_183,w_6_184,w_6_185,w_6_186,w_6_187,w_6_188,w_6_189,w_6_190,w_6_191,w_6_192,w_6_193,w_6_194,w_6_195,w_6_196,w_6_197,w_6_198,w_6_199,w_6_200,w_6_201,w_6_202,w_6_203,w_6_204,w_6_205,w_6_206,w_6_207,w_6_208,w_6_209,w_6_210,w_6_211,w_6_212,w_6_213,w_6_214,w_6_215,w_6_216,w_6_217,w_6_218,w_6_219,w_6_220,w_6_221,w_6_222,w_6_223,w_6_224,w_6_225,w_6_226,w_6_227,w_6_228,w_6_229,w_6_230,w_6_231,w_6_232,w_6_233,w_6_234,w_6_235,w_6_236,w_6_237,w_6_238,w_6_239,w_6_240,w_6_241,w_6_242,w_6_243,w_6_244,w_6_245,w_6_246,w_6_247,w_6_248,w_6_249,w_6_250,w_6_251,w_6_252,w_6_253,w_6_254,w_6_255,w_6_256,w_6_257,w_6_258,w_6_259,w_6_260,w_6_261,w_6_262,w_6_263,w_6_264,w_6_265,w_6_266,w_6_267,w_6_268,w_6_269,w_6_270,w_6_271,w_6_272,w_6_273,w_6_274,w_6_275,w_6_276,w_6_277,w_6_278,w_6_279,w_6_280,w_6_281,w_6_282,w_6_283,w_6_284,w_6_285,w_6_286,w_6_287,w_6_288,w_6_289,w_6_290,w_6_291,w_6_292,w_6_293,w_6_294,w_6_295,w_6_296,w_6_297,w_6_298,w_6_299,w_6_300,w_6_301,w_6_302,w_6_303,w_6_304,w_6_305,w_6_306,w_6_307,w_6_308,w_6_309,w_6_310,w_6_311,w_6_312,w_6_313,w_6_314,w_6_315,w_6_316,w_6_317,w_6_318,w_6_319,w_6_320,w_6_321,w_6_322,w_6_323,w_6_324,w_6_325,w_6_326,w_6_327,w_6_328,w_6_329,w_6_330,w_6_331,w_6_332,w_6_333,w_6_334,w_6_335,w_6_336,w_6_337,w_6_338,w_6_339,w_6_340,w_6_341,w_6_342,w_6_343,w_6_344,w_6_345,w_6_346,w_6_347,w_6_348,w_6_349,w_6_350,w_6_351,w_6_352,w_6_353,w_6_354,w_6_355,w_6_356,w_6_357,w_6_358,w_6_359,w_6_360,w_6_361,w_6_362,w_6_363,w_6_364,w_6_365,w_6_366,w_6_367,w_6_368,w_6_369,w_6_370,w_6_371,w_6_372,w_6_373,w_6_374,w_6_375,w_6_376,w_6_377,w_6_378,w_6_379,w_6_380,w_6_381,w_6_382,w_6_383,w_6_384,w_6_385,w_6_386,w_6_387,w_6_388,w_6_389,w_6_390,w_6_391,w_6_392,w_6_393,w_6_394,w_6_395,w_6_396,w_6_397,w_6_398,w_6_399,w_6_400,w_6_401,w_6_402,w_6_403,w_6_404,w_6_405,w_6_406,w_6_407,w_6_408,w_6_409,w_6_410,w_6_411,w_6_412,w_6_413,w_6_414,w_6_415,w_6_416,w_6_417,w_6_418,w_6_419,w_6_420,w_6_421,w_6_422,w_6_423,w_6_424,w_6_425,w_6_426,w_6_427,w_6_428,w_6_429,w_6_430,w_6_431,w_6_432,w_6_433,w_6_434,w_6_435,w_6_436,w_6_437,w_6_438,w_6_439,w_6_440,w_6_441,w_6_442,w_6_443,w_6_444,w_6_445,w_6_446,w_6_447,w_6_448,w_6_449,w_6_450,w_6_451,w_6_452,w_6_453,w_6_454,w_6_455,w_6_456,w_6_457,w_6_458,w_6_459,w_6_460,w_6_461,w_6_462,w_6_463,w_6_464,w_6_465,w_6_466,w_6_467,w_6_468,w_6_469,w_6_470,w_6_471,w_6_472,w_6_473,w_6_474,w_6_475,w_6_476,w_6_477,w_6_478,w_6_479,w_6_480,w_6_481,w_6_482,w_6_483,w_6_484,w_6_485,w_6_486,w_6_487,w_6_488,w_6_489,w_6_490,w_6_491,w_6_492,w_6_493,w_6_494,w_6_495,w_6_496,w_6_497,w_6_498,w_6_499,w_6_500,w_6_501,w_6_502,w_6_503,w_6_504,w_6_505,w_6_506,w_6_507,w_6_508,w_6_509,w_6_510,w_6_511,w_6_512,w_6_513,w_6_514,w_6_515,w_6_516,w_6_517,w_6_518,w_6_519,w_6_520,w_6_521,w_6_522,w_6_523,w_6_524,w_6_525,w_6_526,w_6_527,w_6_528,w_6_529,w_6_530,w_6_531,w_6_532,w_6_533,w_6_534,w_6_535,w_6_536,w_6_537,w_6_538,w_6_539,w_6_540,w_6_541,w_6_542,w_6_543,w_6_544,w_6_545,w_6_546,w_6_547,w_6_548,w_6_549,w_6_550,w_6_551,w_6_552,w_6_553,w_6_554,w_6_555,w_6_556,w_6_557,w_6_558,w_6_559,w_6_560,w_6_561,w_6_562,w_6_563,w_6_564,w_6_565,w_6_566,w_6_567,w_6_568,w_6_569,w_6_570,w_6_571,w_6_572,w_6_573,w_6_574,w_6_575,w_6_576,w_6_577,w_6_578,w_6_579,w_6_580,w_6_581,w_6_582,w_6_583,w_6_584,w_6_585,w_6_586,w_6_587,w_6_588,w_6_589,w_6_590,w_6_591,w_6_592,w_6_593,w_6_594,w_6_595,w_6_596,w_6_597,w_6_598,w_6_599,w_6_600,w_6_601,w_6_602,w_6_603,w_6_604,w_6_605,w_6_606,w_6_607,w_6_608,w_6_609,w_6_610,w_6_611,w_6_612,w_6_613,w_6_614,w_6_615,w_6_616,w_6_617,w_6_618,w_6_619,w_6_620,w_6_621,w_6_622,w_6_623,w_6_624,w_6_625,w_6_626,w_6_627,w_6_628,w_6_629,w_6_630,w_6_631,w_6_632,w_6_633,w_6_634,w_6_635,w_6_636,w_6_637,w_6_638,w_6_639,w_6_640,w_6_641,w_6_642,w_6_643,w_6_644,w_6_645,w_6_646,w_6_647,w_6_648,w_6_649,w_6_650,w_6_651,w_6_652,w_6_653,w_6_654,w_6_655,w_6_656,w_6_657,w_6_658,w_6_659,w_6_660,w_6_661,w_6_662,w_6_663,w_6_664,w_6_665,w_6_666,w_6_667,w_6_668,w_6_669,w_6_670,w_6_671,w_6_672,w_6_673,w_6_674,w_6_675,w_6_676,w_6_677,w_6_678,w_6_679,w_6_680,w_6_681,w_6_682,w_6_683,w_6_684,w_6_685,w_6_686,w_6_687,w_6_688,w_6_689,w_6_690,w_6_691,w_6_692,w_6_693,w_6_694,w_6_695,w_6_696,w_6_697,w_6_698,w_6_699,w_6_700,w_6_701,w_6_702,w_6_703,w_6_704,w_6_705,w_6_706,w_6_707,w_6_708,w_6_709,w_6_710,w_6_711,w_6_712,w_6_713,w_6_714,w_6_715,w_6_716,w_6_717,w_6_718,w_6_719,w_6_720,w_6_721,w_6_722,w_6_723,w_6_724,w_6_725,w_6_726,w_6_727,w_6_728,w_6_729,w_6_730,w_6_731,w_6_732,w_6_733,w_6_734,w_6_735,w_6_736,w_6_737,w_6_738,w_6_739,w_6_740,w_6_741,w_6_742,w_6_743,w_6_744,w_6_745,w_6_746,w_6_747,w_6_748,w_6_749,w_6_750,w_6_751,w_6_752,w_6_753,w_6_754,w_6_755,w_6_756,w_6_757,w_6_758,w_6_759,w_6_760,w_6_761,w_6_762,w_6_763,w_6_764,w_6_765,w_6_766,w_6_767,w_6_768,w_6_769,w_6_770,w_6_771,w_6_772,w_6_773,w_6_774,w_6_775,w_6_776,w_6_777,w_6_778,w_6_779,w_6_780,w_6_781,w_6_782,w_6_783,w_6_784,
w_7_0,w_7_1,w_7_2,w_7_3,w_7_4,w_7_5,w_7_6,w_7_7,w_7_8,w_7_9,w_7_10,w_7_11,w_7_12,w_7_13,w_7_14,w_7_15,w_7_16,w_7_17,w_7_18,w_7_19,w_7_20,w_7_21,w_7_22,w_7_23,w_7_24,w_7_25,w_7_26,w_7_27,w_7_28,w_7_29,w_7_30,w_7_31,w_7_32,w_7_33,w_7_34,w_7_35,w_7_36,w_7_37,w_7_38,w_7_39,w_7_40,w_7_41,w_7_42,w_7_43,w_7_44,w_7_45,w_7_46,w_7_47,w_7_48,w_7_49,w_7_50,w_7_51,w_7_52,w_7_53,w_7_54,w_7_55,w_7_56,w_7_57,w_7_58,w_7_59,w_7_60,w_7_61,w_7_62,w_7_63,w_7_64,w_7_65,w_7_66,w_7_67,w_7_68,w_7_69,w_7_70,w_7_71,w_7_72,w_7_73,w_7_74,w_7_75,w_7_76,w_7_77,w_7_78,w_7_79,w_7_80,w_7_81,w_7_82,w_7_83,w_7_84,w_7_85,w_7_86,w_7_87,w_7_88,w_7_89,w_7_90,w_7_91,w_7_92,w_7_93,w_7_94,w_7_95,w_7_96,w_7_97,w_7_98,w_7_99,w_7_100,w_7_101,w_7_102,w_7_103,w_7_104,w_7_105,w_7_106,w_7_107,w_7_108,w_7_109,w_7_110,w_7_111,w_7_112,w_7_113,w_7_114,w_7_115,w_7_116,w_7_117,w_7_118,w_7_119,w_7_120,w_7_121,w_7_122,w_7_123,w_7_124,w_7_125,w_7_126,w_7_127,w_7_128,w_7_129,w_7_130,w_7_131,w_7_132,w_7_133,w_7_134,w_7_135,w_7_136,w_7_137,w_7_138,w_7_139,w_7_140,w_7_141,w_7_142,w_7_143,w_7_144,w_7_145,w_7_146,w_7_147,w_7_148,w_7_149,w_7_150,w_7_151,w_7_152,w_7_153,w_7_154,w_7_155,w_7_156,w_7_157,w_7_158,w_7_159,w_7_160,w_7_161,w_7_162,w_7_163,w_7_164,w_7_165,w_7_166,w_7_167,w_7_168,w_7_169,w_7_170,w_7_171,w_7_172,w_7_173,w_7_174,w_7_175,w_7_176,w_7_177,w_7_178,w_7_179,w_7_180,w_7_181,w_7_182,w_7_183,w_7_184,w_7_185,w_7_186,w_7_187,w_7_188,w_7_189,w_7_190,w_7_191,w_7_192,w_7_193,w_7_194,w_7_195,w_7_196,w_7_197,w_7_198,w_7_199,w_7_200,w_7_201,w_7_202,w_7_203,w_7_204,w_7_205,w_7_206,w_7_207,w_7_208,w_7_209,w_7_210,w_7_211,w_7_212,w_7_213,w_7_214,w_7_215,w_7_216,w_7_217,w_7_218,w_7_219,w_7_220,w_7_221,w_7_222,w_7_223,w_7_224,w_7_225,w_7_226,w_7_227,w_7_228,w_7_229,w_7_230,w_7_231,w_7_232,w_7_233,w_7_234,w_7_235,w_7_236,w_7_237,w_7_238,w_7_239,w_7_240,w_7_241,w_7_242,w_7_243,w_7_244,w_7_245,w_7_246,w_7_247,w_7_248,w_7_249,w_7_250,w_7_251,w_7_252,w_7_253,w_7_254,w_7_255,w_7_256,w_7_257,w_7_258,w_7_259,w_7_260,w_7_261,w_7_262,w_7_263,w_7_264,w_7_265,w_7_266,w_7_267,w_7_268,w_7_269,w_7_270,w_7_271,w_7_272,w_7_273,w_7_274,w_7_275,w_7_276,w_7_277,w_7_278,w_7_279,w_7_280,w_7_281,w_7_282,w_7_283,w_7_284,w_7_285,w_7_286,w_7_287,w_7_288,w_7_289,w_7_290,w_7_291,w_7_292,w_7_293,w_7_294,w_7_295,w_7_296,w_7_297,w_7_298,w_7_299,w_7_300,w_7_301,w_7_302,w_7_303,w_7_304,w_7_305,w_7_306,w_7_307,w_7_308,w_7_309,w_7_310,w_7_311,w_7_312,w_7_313,w_7_314,w_7_315,w_7_316,w_7_317,w_7_318,w_7_319,w_7_320,w_7_321,w_7_322,w_7_323,w_7_324,w_7_325,w_7_326,w_7_327,w_7_328,w_7_329,w_7_330,w_7_331,w_7_332,w_7_333,w_7_334,w_7_335,w_7_336,w_7_337,w_7_338,w_7_339,w_7_340,w_7_341,w_7_342,w_7_343,w_7_344,w_7_345,w_7_346,w_7_347,w_7_348,w_7_349,w_7_350,w_7_351,w_7_352,w_7_353,w_7_354,w_7_355,w_7_356,w_7_357,w_7_358,w_7_359,w_7_360,w_7_361,w_7_362,w_7_363,w_7_364,w_7_365,w_7_366,w_7_367,w_7_368,w_7_369,w_7_370,w_7_371,w_7_372,w_7_373,w_7_374,w_7_375,w_7_376,w_7_377,w_7_378,w_7_379,w_7_380,w_7_381,w_7_382,w_7_383,w_7_384,w_7_385,w_7_386,w_7_387,w_7_388,w_7_389,w_7_390,w_7_391,w_7_392,w_7_393,w_7_394,w_7_395,w_7_396,w_7_397,w_7_398,w_7_399,w_7_400,w_7_401,w_7_402,w_7_403,w_7_404,w_7_405,w_7_406,w_7_407,w_7_408,w_7_409,w_7_410,w_7_411,w_7_412,w_7_413,w_7_414,w_7_415,w_7_416,w_7_417,w_7_418,w_7_419,w_7_420,w_7_421,w_7_422,w_7_423,w_7_424,w_7_425,w_7_426,w_7_427,w_7_428,w_7_429,w_7_430,w_7_431,w_7_432,w_7_433,w_7_434,w_7_435,w_7_436,w_7_437,w_7_438,w_7_439,w_7_440,w_7_441,w_7_442,w_7_443,w_7_444,w_7_445,w_7_446,w_7_447,w_7_448,w_7_449,w_7_450,w_7_451,w_7_452,w_7_453,w_7_454,w_7_455,w_7_456,w_7_457,w_7_458,w_7_459,w_7_460,w_7_461,w_7_462,w_7_463,w_7_464,w_7_465,w_7_466,w_7_467,w_7_468,w_7_469,w_7_470,w_7_471,w_7_472,w_7_473,w_7_474,w_7_475,w_7_476,w_7_477,w_7_478,w_7_479,w_7_480,w_7_481,w_7_482,w_7_483,w_7_484,w_7_485,w_7_486,w_7_487,w_7_488,w_7_489,w_7_490,w_7_491,w_7_492,w_7_493,w_7_494,w_7_495,w_7_496,w_7_497,w_7_498,w_7_499,w_7_500,w_7_501,w_7_502,w_7_503,w_7_504,w_7_505,w_7_506,w_7_507,w_7_508,w_7_509,w_7_510,w_7_511,w_7_512,w_7_513,w_7_514,w_7_515,w_7_516,w_7_517,w_7_518,w_7_519,w_7_520,w_7_521,w_7_522,w_7_523,w_7_524,w_7_525,w_7_526,w_7_527,w_7_528,w_7_529,w_7_530,w_7_531,w_7_532,w_7_533,w_7_534,w_7_535,w_7_536,w_7_537,w_7_538,w_7_539,w_7_540,w_7_541,w_7_542,w_7_543,w_7_544,w_7_545,w_7_546,w_7_547,w_7_548,w_7_549,w_7_550,w_7_551,w_7_552,w_7_553,w_7_554,w_7_555,w_7_556,w_7_557,w_7_558,w_7_559,w_7_560,w_7_561,w_7_562,w_7_563,w_7_564,w_7_565,w_7_566,w_7_567,w_7_568,w_7_569,w_7_570,w_7_571,w_7_572,w_7_573,w_7_574,w_7_575,w_7_576,w_7_577,w_7_578,w_7_579,w_7_580,w_7_581,w_7_582,w_7_583,w_7_584,w_7_585,w_7_586,w_7_587,w_7_588,w_7_589,w_7_590,w_7_591,w_7_592,w_7_593,w_7_594,w_7_595,w_7_596,w_7_597,w_7_598,w_7_599,w_7_600,w_7_601,w_7_602,w_7_603,w_7_604,w_7_605,w_7_606,w_7_607,w_7_608,w_7_609,w_7_610,w_7_611,w_7_612,w_7_613,w_7_614,w_7_615,w_7_616,w_7_617,w_7_618,w_7_619,w_7_620,w_7_621,w_7_622,w_7_623,w_7_624,w_7_625,w_7_626,w_7_627,w_7_628,w_7_629,w_7_630,w_7_631,w_7_632,w_7_633,w_7_634,w_7_635,w_7_636,w_7_637,w_7_638,w_7_639,w_7_640,w_7_641,w_7_642,w_7_643,w_7_644,w_7_645,w_7_646,w_7_647,w_7_648,w_7_649,w_7_650,w_7_651,w_7_652,w_7_653,w_7_654,w_7_655,w_7_656,w_7_657,w_7_658,w_7_659,w_7_660,w_7_661,w_7_662,w_7_663,w_7_664,w_7_665,w_7_666,w_7_667,w_7_668,w_7_669,w_7_670,w_7_671,w_7_672,w_7_673,w_7_674,w_7_675,w_7_676,w_7_677,w_7_678,w_7_679,w_7_680,w_7_681,w_7_682,w_7_683,w_7_684,w_7_685,w_7_686,w_7_687,w_7_688,w_7_689,w_7_690,w_7_691,w_7_692,w_7_693,w_7_694,w_7_695,w_7_696,w_7_697,w_7_698,w_7_699,w_7_700,w_7_701,w_7_702,w_7_703,w_7_704,w_7_705,w_7_706,w_7_707,w_7_708,w_7_709,w_7_710,w_7_711,w_7_712,w_7_713,w_7_714,w_7_715,w_7_716,w_7_717,w_7_718,w_7_719,w_7_720,w_7_721,w_7_722,w_7_723,w_7_724,w_7_725,w_7_726,w_7_727,w_7_728,w_7_729,w_7_730,w_7_731,w_7_732,w_7_733,w_7_734,w_7_735,w_7_736,w_7_737,w_7_738,w_7_739,w_7_740,w_7_741,w_7_742,w_7_743,w_7_744,w_7_745,w_7_746,w_7_747,w_7_748,w_7_749,w_7_750,w_7_751,w_7_752,w_7_753,w_7_754,w_7_755,w_7_756,w_7_757,w_7_758,w_7_759,w_7_760,w_7_761,w_7_762,w_7_763,w_7_764,w_7_765,w_7_766,w_7_767,w_7_768,w_7_769,w_7_770,w_7_771,w_7_772,w_7_773,w_7_774,w_7_775,w_7_776,w_7_777,w_7_778,w_7_779,w_7_780,w_7_781,w_7_782,w_7_783,w_7_784,
w_8_0,w_8_1,w_8_2,w_8_3,w_8_4,w_8_5,w_8_6,w_8_7,w_8_8,w_8_9,w_8_10,w_8_11,w_8_12,w_8_13,w_8_14,w_8_15,w_8_16,w_8_17,w_8_18,w_8_19,w_8_20,w_8_21,w_8_22,w_8_23,w_8_24,w_8_25,w_8_26,w_8_27,w_8_28,w_8_29,w_8_30,w_8_31,w_8_32,w_8_33,w_8_34,w_8_35,w_8_36,w_8_37,w_8_38,w_8_39,w_8_40,w_8_41,w_8_42,w_8_43,w_8_44,w_8_45,w_8_46,w_8_47,w_8_48,w_8_49,w_8_50,w_8_51,w_8_52,w_8_53,w_8_54,w_8_55,w_8_56,w_8_57,w_8_58,w_8_59,w_8_60,w_8_61,w_8_62,w_8_63,w_8_64,w_8_65,w_8_66,w_8_67,w_8_68,w_8_69,w_8_70,w_8_71,w_8_72,w_8_73,w_8_74,w_8_75,w_8_76,w_8_77,w_8_78,w_8_79,w_8_80,w_8_81,w_8_82,w_8_83,w_8_84,w_8_85,w_8_86,w_8_87,w_8_88,w_8_89,w_8_90,w_8_91,w_8_92,w_8_93,w_8_94,w_8_95,w_8_96,w_8_97,w_8_98,w_8_99,w_8_100,w_8_101,w_8_102,w_8_103,w_8_104,w_8_105,w_8_106,w_8_107,w_8_108,w_8_109,w_8_110,w_8_111,w_8_112,w_8_113,w_8_114,w_8_115,w_8_116,w_8_117,w_8_118,w_8_119,w_8_120,w_8_121,w_8_122,w_8_123,w_8_124,w_8_125,w_8_126,w_8_127,w_8_128,w_8_129,w_8_130,w_8_131,w_8_132,w_8_133,w_8_134,w_8_135,w_8_136,w_8_137,w_8_138,w_8_139,w_8_140,w_8_141,w_8_142,w_8_143,w_8_144,w_8_145,w_8_146,w_8_147,w_8_148,w_8_149,w_8_150,w_8_151,w_8_152,w_8_153,w_8_154,w_8_155,w_8_156,w_8_157,w_8_158,w_8_159,w_8_160,w_8_161,w_8_162,w_8_163,w_8_164,w_8_165,w_8_166,w_8_167,w_8_168,w_8_169,w_8_170,w_8_171,w_8_172,w_8_173,w_8_174,w_8_175,w_8_176,w_8_177,w_8_178,w_8_179,w_8_180,w_8_181,w_8_182,w_8_183,w_8_184,w_8_185,w_8_186,w_8_187,w_8_188,w_8_189,w_8_190,w_8_191,w_8_192,w_8_193,w_8_194,w_8_195,w_8_196,w_8_197,w_8_198,w_8_199,w_8_200,w_8_201,w_8_202,w_8_203,w_8_204,w_8_205,w_8_206,w_8_207,w_8_208,w_8_209,w_8_210,w_8_211,w_8_212,w_8_213,w_8_214,w_8_215,w_8_216,w_8_217,w_8_218,w_8_219,w_8_220,w_8_221,w_8_222,w_8_223,w_8_224,w_8_225,w_8_226,w_8_227,w_8_228,w_8_229,w_8_230,w_8_231,w_8_232,w_8_233,w_8_234,w_8_235,w_8_236,w_8_237,w_8_238,w_8_239,w_8_240,w_8_241,w_8_242,w_8_243,w_8_244,w_8_245,w_8_246,w_8_247,w_8_248,w_8_249,w_8_250,w_8_251,w_8_252,w_8_253,w_8_254,w_8_255,w_8_256,w_8_257,w_8_258,w_8_259,w_8_260,w_8_261,w_8_262,w_8_263,w_8_264,w_8_265,w_8_266,w_8_267,w_8_268,w_8_269,w_8_270,w_8_271,w_8_272,w_8_273,w_8_274,w_8_275,w_8_276,w_8_277,w_8_278,w_8_279,w_8_280,w_8_281,w_8_282,w_8_283,w_8_284,w_8_285,w_8_286,w_8_287,w_8_288,w_8_289,w_8_290,w_8_291,w_8_292,w_8_293,w_8_294,w_8_295,w_8_296,w_8_297,w_8_298,w_8_299,w_8_300,w_8_301,w_8_302,w_8_303,w_8_304,w_8_305,w_8_306,w_8_307,w_8_308,w_8_309,w_8_310,w_8_311,w_8_312,w_8_313,w_8_314,w_8_315,w_8_316,w_8_317,w_8_318,w_8_319,w_8_320,w_8_321,w_8_322,w_8_323,w_8_324,w_8_325,w_8_326,w_8_327,w_8_328,w_8_329,w_8_330,w_8_331,w_8_332,w_8_333,w_8_334,w_8_335,w_8_336,w_8_337,w_8_338,w_8_339,w_8_340,w_8_341,w_8_342,w_8_343,w_8_344,w_8_345,w_8_346,w_8_347,w_8_348,w_8_349,w_8_350,w_8_351,w_8_352,w_8_353,w_8_354,w_8_355,w_8_356,w_8_357,w_8_358,w_8_359,w_8_360,w_8_361,w_8_362,w_8_363,w_8_364,w_8_365,w_8_366,w_8_367,w_8_368,w_8_369,w_8_370,w_8_371,w_8_372,w_8_373,w_8_374,w_8_375,w_8_376,w_8_377,w_8_378,w_8_379,w_8_380,w_8_381,w_8_382,w_8_383,w_8_384,w_8_385,w_8_386,w_8_387,w_8_388,w_8_389,w_8_390,w_8_391,w_8_392,w_8_393,w_8_394,w_8_395,w_8_396,w_8_397,w_8_398,w_8_399,w_8_400,w_8_401,w_8_402,w_8_403,w_8_404,w_8_405,w_8_406,w_8_407,w_8_408,w_8_409,w_8_410,w_8_411,w_8_412,w_8_413,w_8_414,w_8_415,w_8_416,w_8_417,w_8_418,w_8_419,w_8_420,w_8_421,w_8_422,w_8_423,w_8_424,w_8_425,w_8_426,w_8_427,w_8_428,w_8_429,w_8_430,w_8_431,w_8_432,w_8_433,w_8_434,w_8_435,w_8_436,w_8_437,w_8_438,w_8_439,w_8_440,w_8_441,w_8_442,w_8_443,w_8_444,w_8_445,w_8_446,w_8_447,w_8_448,w_8_449,w_8_450,w_8_451,w_8_452,w_8_453,w_8_454,w_8_455,w_8_456,w_8_457,w_8_458,w_8_459,w_8_460,w_8_461,w_8_462,w_8_463,w_8_464,w_8_465,w_8_466,w_8_467,w_8_468,w_8_469,w_8_470,w_8_471,w_8_472,w_8_473,w_8_474,w_8_475,w_8_476,w_8_477,w_8_478,w_8_479,w_8_480,w_8_481,w_8_482,w_8_483,w_8_484,w_8_485,w_8_486,w_8_487,w_8_488,w_8_489,w_8_490,w_8_491,w_8_492,w_8_493,w_8_494,w_8_495,w_8_496,w_8_497,w_8_498,w_8_499,w_8_500,w_8_501,w_8_502,w_8_503,w_8_504,w_8_505,w_8_506,w_8_507,w_8_508,w_8_509,w_8_510,w_8_511,w_8_512,w_8_513,w_8_514,w_8_515,w_8_516,w_8_517,w_8_518,w_8_519,w_8_520,w_8_521,w_8_522,w_8_523,w_8_524,w_8_525,w_8_526,w_8_527,w_8_528,w_8_529,w_8_530,w_8_531,w_8_532,w_8_533,w_8_534,w_8_535,w_8_536,w_8_537,w_8_538,w_8_539,w_8_540,w_8_541,w_8_542,w_8_543,w_8_544,w_8_545,w_8_546,w_8_547,w_8_548,w_8_549,w_8_550,w_8_551,w_8_552,w_8_553,w_8_554,w_8_555,w_8_556,w_8_557,w_8_558,w_8_559,w_8_560,w_8_561,w_8_562,w_8_563,w_8_564,w_8_565,w_8_566,w_8_567,w_8_568,w_8_569,w_8_570,w_8_571,w_8_572,w_8_573,w_8_574,w_8_575,w_8_576,w_8_577,w_8_578,w_8_579,w_8_580,w_8_581,w_8_582,w_8_583,w_8_584,w_8_585,w_8_586,w_8_587,w_8_588,w_8_589,w_8_590,w_8_591,w_8_592,w_8_593,w_8_594,w_8_595,w_8_596,w_8_597,w_8_598,w_8_599,w_8_600,w_8_601,w_8_602,w_8_603,w_8_604,w_8_605,w_8_606,w_8_607,w_8_608,w_8_609,w_8_610,w_8_611,w_8_612,w_8_613,w_8_614,w_8_615,w_8_616,w_8_617,w_8_618,w_8_619,w_8_620,w_8_621,w_8_622,w_8_623,w_8_624,w_8_625,w_8_626,w_8_627,w_8_628,w_8_629,w_8_630,w_8_631,w_8_632,w_8_633,w_8_634,w_8_635,w_8_636,w_8_637,w_8_638,w_8_639,w_8_640,w_8_641,w_8_642,w_8_643,w_8_644,w_8_645,w_8_646,w_8_647,w_8_648,w_8_649,w_8_650,w_8_651,w_8_652,w_8_653,w_8_654,w_8_655,w_8_656,w_8_657,w_8_658,w_8_659,w_8_660,w_8_661,w_8_662,w_8_663,w_8_664,w_8_665,w_8_666,w_8_667,w_8_668,w_8_669,w_8_670,w_8_671,w_8_672,w_8_673,w_8_674,w_8_675,w_8_676,w_8_677,w_8_678,w_8_679,w_8_680,w_8_681,w_8_682,w_8_683,w_8_684,w_8_685,w_8_686,w_8_687,w_8_688,w_8_689,w_8_690,w_8_691,w_8_692,w_8_693,w_8_694,w_8_695,w_8_696,w_8_697,w_8_698,w_8_699,w_8_700,w_8_701,w_8_702,w_8_703,w_8_704,w_8_705,w_8_706,w_8_707,w_8_708,w_8_709,w_8_710,w_8_711,w_8_712,w_8_713,w_8_714,w_8_715,w_8_716,w_8_717,w_8_718,w_8_719,w_8_720,w_8_721,w_8_722,w_8_723,w_8_724,w_8_725,w_8_726,w_8_727,w_8_728,w_8_729,w_8_730,w_8_731,w_8_732,w_8_733,w_8_734,w_8_735,w_8_736,w_8_737,w_8_738,w_8_739,w_8_740,w_8_741,w_8_742,w_8_743,w_8_744,w_8_745,w_8_746,w_8_747,w_8_748,w_8_749,w_8_750,w_8_751,w_8_752,w_8_753,w_8_754,w_8_755,w_8_756,w_8_757,w_8_758,w_8_759,w_8_760,w_8_761,w_8_762,w_8_763,w_8_764,w_8_765,w_8_766,w_8_767,w_8_768,w_8_769,w_8_770,w_8_771,w_8_772,w_8_773,w_8_774,w_8_775,w_8_776,w_8_777,w_8_778,w_8_779,w_8_780,w_8_781,w_8_782,w_8_783,w_8_784,
w_9_0,w_9_1,w_9_2,w_9_3,w_9_4,w_9_5,w_9_6,w_9_7,w_9_8,w_9_9,w_9_10,w_9_11,w_9_12,w_9_13,w_9_14,w_9_15,w_9_16,w_9_17,w_9_18,w_9_19,w_9_20,w_9_21,w_9_22,w_9_23,w_9_24,w_9_25,w_9_26,w_9_27,w_9_28,w_9_29,w_9_30,w_9_31,w_9_32,w_9_33,w_9_34,w_9_35,w_9_36,w_9_37,w_9_38,w_9_39,w_9_40,w_9_41,w_9_42,w_9_43,w_9_44,w_9_45,w_9_46,w_9_47,w_9_48,w_9_49,w_9_50,w_9_51,w_9_52,w_9_53,w_9_54,w_9_55,w_9_56,w_9_57,w_9_58,w_9_59,w_9_60,w_9_61,w_9_62,w_9_63,w_9_64,w_9_65,w_9_66,w_9_67,w_9_68,w_9_69,w_9_70,w_9_71,w_9_72,w_9_73,w_9_74,w_9_75,w_9_76,w_9_77,w_9_78,w_9_79,w_9_80,w_9_81,w_9_82,w_9_83,w_9_84,w_9_85,w_9_86,w_9_87,w_9_88,w_9_89,w_9_90,w_9_91,w_9_92,w_9_93,w_9_94,w_9_95,w_9_96,w_9_97,w_9_98,w_9_99,w_9_100,w_9_101,w_9_102,w_9_103,w_9_104,w_9_105,w_9_106,w_9_107,w_9_108,w_9_109,w_9_110,w_9_111,w_9_112,w_9_113,w_9_114,w_9_115,w_9_116,w_9_117,w_9_118,w_9_119,w_9_120,w_9_121,w_9_122,w_9_123,w_9_124,w_9_125,w_9_126,w_9_127,w_9_128,w_9_129,w_9_130,w_9_131,w_9_132,w_9_133,w_9_134,w_9_135,w_9_136,w_9_137,w_9_138,w_9_139,w_9_140,w_9_141,w_9_142,w_9_143,w_9_144,w_9_145,w_9_146,w_9_147,w_9_148,w_9_149,w_9_150,w_9_151,w_9_152,w_9_153,w_9_154,w_9_155,w_9_156,w_9_157,w_9_158,w_9_159,w_9_160,w_9_161,w_9_162,w_9_163,w_9_164,w_9_165,w_9_166,w_9_167,w_9_168,w_9_169,w_9_170,w_9_171,w_9_172,w_9_173,w_9_174,w_9_175,w_9_176,w_9_177,w_9_178,w_9_179,w_9_180,w_9_181,w_9_182,w_9_183,w_9_184,w_9_185,w_9_186,w_9_187,w_9_188,w_9_189,w_9_190,w_9_191,w_9_192,w_9_193,w_9_194,w_9_195,w_9_196,w_9_197,w_9_198,w_9_199,w_9_200,w_9_201,w_9_202,w_9_203,w_9_204,w_9_205,w_9_206,w_9_207,w_9_208,w_9_209,w_9_210,w_9_211,w_9_212,w_9_213,w_9_214,w_9_215,w_9_216,w_9_217,w_9_218,w_9_219,w_9_220,w_9_221,w_9_222,w_9_223,w_9_224,w_9_225,w_9_226,w_9_227,w_9_228,w_9_229,w_9_230,w_9_231,w_9_232,w_9_233,w_9_234,w_9_235,w_9_236,w_9_237,w_9_238,w_9_239,w_9_240,w_9_241,w_9_242,w_9_243,w_9_244,w_9_245,w_9_246,w_9_247,w_9_248,w_9_249,w_9_250,w_9_251,w_9_252,w_9_253,w_9_254,w_9_255,w_9_256,w_9_257,w_9_258,w_9_259,w_9_260,w_9_261,w_9_262,w_9_263,w_9_264,w_9_265,w_9_266,w_9_267,w_9_268,w_9_269,w_9_270,w_9_271,w_9_272,w_9_273,w_9_274,w_9_275,w_9_276,w_9_277,w_9_278,w_9_279,w_9_280,w_9_281,w_9_282,w_9_283,w_9_284,w_9_285,w_9_286,w_9_287,w_9_288,w_9_289,w_9_290,w_9_291,w_9_292,w_9_293,w_9_294,w_9_295,w_9_296,w_9_297,w_9_298,w_9_299,w_9_300,w_9_301,w_9_302,w_9_303,w_9_304,w_9_305,w_9_306,w_9_307,w_9_308,w_9_309,w_9_310,w_9_311,w_9_312,w_9_313,w_9_314,w_9_315,w_9_316,w_9_317,w_9_318,w_9_319,w_9_320,w_9_321,w_9_322,w_9_323,w_9_324,w_9_325,w_9_326,w_9_327,w_9_328,w_9_329,w_9_330,w_9_331,w_9_332,w_9_333,w_9_334,w_9_335,w_9_336,w_9_337,w_9_338,w_9_339,w_9_340,w_9_341,w_9_342,w_9_343,w_9_344,w_9_345,w_9_346,w_9_347,w_9_348,w_9_349,w_9_350,w_9_351,w_9_352,w_9_353,w_9_354,w_9_355,w_9_356,w_9_357,w_9_358,w_9_359,w_9_360,w_9_361,w_9_362,w_9_363,w_9_364,w_9_365,w_9_366,w_9_367,w_9_368,w_9_369,w_9_370,w_9_371,w_9_372,w_9_373,w_9_374,w_9_375,w_9_376,w_9_377,w_9_378,w_9_379,w_9_380,w_9_381,w_9_382,w_9_383,w_9_384,w_9_385,w_9_386,w_9_387,w_9_388,w_9_389,w_9_390,w_9_391,w_9_392,w_9_393,w_9_394,w_9_395,w_9_396,w_9_397,w_9_398,w_9_399,w_9_400,w_9_401,w_9_402,w_9_403,w_9_404,w_9_405,w_9_406,w_9_407,w_9_408,w_9_409,w_9_410,w_9_411,w_9_412,w_9_413,w_9_414,w_9_415,w_9_416,w_9_417,w_9_418,w_9_419,w_9_420,w_9_421,w_9_422,w_9_423,w_9_424,w_9_425,w_9_426,w_9_427,w_9_428,w_9_429,w_9_430,w_9_431,w_9_432,w_9_433,w_9_434,w_9_435,w_9_436,w_9_437,w_9_438,w_9_439,w_9_440,w_9_441,w_9_442,w_9_443,w_9_444,w_9_445,w_9_446,w_9_447,w_9_448,w_9_449,w_9_450,w_9_451,w_9_452,w_9_453,w_9_454,w_9_455,w_9_456,w_9_457,w_9_458,w_9_459,w_9_460,w_9_461,w_9_462,w_9_463,w_9_464,w_9_465,w_9_466,w_9_467,w_9_468,w_9_469,w_9_470,w_9_471,w_9_472,w_9_473,w_9_474,w_9_475,w_9_476,w_9_477,w_9_478,w_9_479,w_9_480,w_9_481,w_9_482,w_9_483,w_9_484,w_9_485,w_9_486,w_9_487,w_9_488,w_9_489,w_9_490,w_9_491,w_9_492,w_9_493,w_9_494,w_9_495,w_9_496,w_9_497,w_9_498,w_9_499,w_9_500,w_9_501,w_9_502,w_9_503,w_9_504,w_9_505,w_9_506,w_9_507,w_9_508,w_9_509,w_9_510,w_9_511,w_9_512,w_9_513,w_9_514,w_9_515,w_9_516,w_9_517,w_9_518,w_9_519,w_9_520,w_9_521,w_9_522,w_9_523,w_9_524,w_9_525,w_9_526,w_9_527,w_9_528,w_9_529,w_9_530,w_9_531,w_9_532,w_9_533,w_9_534,w_9_535,w_9_536,w_9_537,w_9_538,w_9_539,w_9_540,w_9_541,w_9_542,w_9_543,w_9_544,w_9_545,w_9_546,w_9_547,w_9_548,w_9_549,w_9_550,w_9_551,w_9_552,w_9_553,w_9_554,w_9_555,w_9_556,w_9_557,w_9_558,w_9_559,w_9_560,w_9_561,w_9_562,w_9_563,w_9_564,w_9_565,w_9_566,w_9_567,w_9_568,w_9_569,w_9_570,w_9_571,w_9_572,w_9_573,w_9_574,w_9_575,w_9_576,w_9_577,w_9_578,w_9_579,w_9_580,w_9_581,w_9_582,w_9_583,w_9_584,w_9_585,w_9_586,w_9_587,w_9_588,w_9_589,w_9_590,w_9_591,w_9_592,w_9_593,w_9_594,w_9_595,w_9_596,w_9_597,w_9_598,w_9_599,w_9_600,w_9_601,w_9_602,w_9_603,w_9_604,w_9_605,w_9_606,w_9_607,w_9_608,w_9_609,w_9_610,w_9_611,w_9_612,w_9_613,w_9_614,w_9_615,w_9_616,w_9_617,w_9_618,w_9_619,w_9_620,w_9_621,w_9_622,w_9_623,w_9_624,w_9_625,w_9_626,w_9_627,w_9_628,w_9_629,w_9_630,w_9_631,w_9_632,w_9_633,w_9_634,w_9_635,w_9_636,w_9_637,w_9_638,w_9_639,w_9_640,w_9_641,w_9_642,w_9_643,w_9_644,w_9_645,w_9_646,w_9_647,w_9_648,w_9_649,w_9_650,w_9_651,w_9_652,w_9_653,w_9_654,w_9_655,w_9_656,w_9_657,w_9_658,w_9_659,w_9_660,w_9_661,w_9_662,w_9_663,w_9_664,w_9_665,w_9_666,w_9_667,w_9_668,w_9_669,w_9_670,w_9_671,w_9_672,w_9_673,w_9_674,w_9_675,w_9_676,w_9_677,w_9_678,w_9_679,w_9_680,w_9_681,w_9_682,w_9_683,w_9_684,w_9_685,w_9_686,w_9_687,w_9_688,w_9_689,w_9_690,w_9_691,w_9_692,w_9_693,w_9_694,w_9_695,w_9_696,w_9_697,w_9_698,w_9_699,w_9_700,w_9_701,w_9_702,w_9_703,w_9_704,w_9_705,w_9_706,w_9_707,w_9_708,w_9_709,w_9_710,w_9_711,w_9_712,w_9_713,w_9_714,w_9_715,w_9_716,w_9_717,w_9_718,w_9_719,w_9_720,w_9_721,w_9_722,w_9_723,w_9_724,w_9_725,w_9_726,w_9_727,w_9_728,w_9_729,w_9_730,w_9_731,w_9_732,w_9_733,w_9_734,w_9_735,w_9_736,w_9_737,w_9_738,w_9_739,w_9_740,w_9_741,w_9_742,w_9_743,w_9_744,w_9_745,w_9_746,w_9_747,w_9_748,w_9_749,w_9_750,w_9_751,w_9_752,w_9_753,w_9_754,w_9_755,w_9_756,w_9_757,w_9_758,w_9_759,w_9_760,w_9_761,w_9_762,w_9_763,w_9_764,w_9_765,w_9_766,w_9_767,w_9_768,w_9_769,w_9_770,w_9_771,w_9_772,w_9_773,w_9_774,w_9_775,w_9_776,w_9_777,w_9_778,w_9_779,w_9_780,w_9_781,w_9_782,w_9_783,w_9_784;

reg [9:0] px_0,px_1,px_2,px_3,px_4,px_5,px_6,px_7,px_8,px_9,px_10,px_11,px_12,px_13,px_14,px_15,px_16,px_17,px_18,px_19,px_20,px_21,px_22,px_23,px_24,px_25,px_26,px_27,px_28,px_29,px_30,px_31,px_32,px_33,px_34,px_35,px_36,px_37,px_38,px_39,px_40,px_41,px_42,px_43,px_44,px_45,px_46,px_47,px_48,px_49,px_50,px_51,px_52,px_53,px_54,px_55,px_56,px_57,px_58,px_59,px_60,px_61,px_62,px_63,px_64,px_65,px_66,px_67,px_68,px_69,px_70,px_71,px_72,px_73,px_74,px_75,px_76,px_77,px_78,px_79,px_80,px_81,px_82,px_83,px_84,px_85,px_86,px_87,px_88,px_89,px_90,px_91,px_92,px_93,px_94,px_95,px_96,px_97,px_98,px_99,px_100,px_101,px_102,px_103,px_104,px_105,px_106,px_107,px_108,px_109,px_110,px_111,px_112,px_113,px_114,px_115,px_116,px_117,px_118,px_119,px_120,px_121,px_122,px_123,px_124,px_125,px_126,px_127,px_128,px_129,px_130,px_131,px_132,px_133,px_134,px_135,px_136,px_137,px_138,px_139,px_140,px_141,px_142,px_143,px_144,px_145,px_146,px_147,px_148,px_149,px_150,px_151,px_152,px_153,px_154,px_155,px_156,px_157,px_158,px_159,px_160,px_161,px_162,px_163,px_164,px_165,px_166,px_167,px_168,px_169,px_170,px_171,px_172,px_173,px_174,px_175,px_176,px_177,px_178,px_179,px_180,px_181,px_182,px_183,px_184,px_185,px_186,px_187,px_188,px_189,px_190,px_191,px_192,px_193,px_194,px_195,px_196,px_197,px_198,px_199,px_200,px_201,px_202,px_203,px_204,px_205,px_206,px_207,px_208,px_209,px_210,px_211,px_212,px_213,px_214,px_215,px_216,px_217,px_218,px_219,px_220,px_221,px_222,px_223,px_224,px_225,px_226,px_227,px_228,px_229,px_230,px_231,px_232,px_233,px_234,px_235,px_236,px_237,px_238,px_239,px_240,px_241,px_242,px_243,px_244,px_245,px_246,px_247,px_248,px_249,px_250,px_251,px_252,px_253,px_254,px_255,px_256,px_257,px_258,px_259,px_260,px_261,px_262,px_263,px_264,px_265,px_266,px_267,px_268,px_269,px_270,px_271,px_272,px_273,px_274,px_275,px_276,px_277,px_278,px_279,px_280,px_281,px_282,px_283,px_284,px_285,px_286,px_287,px_288,px_289,px_290,px_291,px_292,px_293,px_294,px_295,px_296,px_297,px_298,px_299,px_300,px_301,px_302,px_303,px_304,px_305,px_306,px_307,px_308,px_309,px_310,px_311,px_312,px_313,px_314,px_315,px_316,px_317,px_318,px_319,px_320,px_321,px_322,px_323,px_324,px_325,px_326,px_327,px_328,px_329,px_330,px_331,px_332,px_333,px_334,px_335,px_336,px_337,px_338,px_339,px_340,px_341,px_342,px_343,px_344,px_345,px_346,px_347,px_348,px_349,px_350,px_351,px_352,px_353,px_354,px_355,px_356,px_357,px_358,px_359,px_360,px_361,px_362,px_363,px_364,px_365,px_366,px_367,px_368,px_369,px_370,px_371,px_372,px_373,px_374,px_375,px_376,px_377,px_378,px_379,px_380,px_381,px_382,px_383,px_384,px_385,px_386,px_387,px_388,px_389,px_390,px_391,px_392,px_393,px_394,px_395,px_396,px_397,px_398,px_399,px_400,px_401,px_402,px_403,px_404,px_405,px_406,px_407,px_408,px_409,px_410,px_411,px_412,px_413,px_414,px_415,px_416,px_417,px_418,px_419,px_420,px_421,px_422,px_423,px_424,px_425,px_426,px_427,px_428,px_429,px_430,px_431,px_432,px_433,px_434,px_435,px_436,px_437,px_438,px_439,px_440,px_441,px_442,px_443,px_444,px_445,px_446,px_447,px_448,px_449,px_450,px_451,px_452,px_453,px_454,px_455,px_456,px_457,px_458,px_459,px_460,px_461,px_462,px_463,px_464,px_465,px_466,px_467,px_468,px_469,px_470,px_471,px_472,px_473,px_474,px_475,px_476,px_477,px_478,px_479,px_480,px_481,px_482,px_483,px_484,px_485,px_486,px_487,px_488,px_489,px_490,px_491,px_492,px_493,px_494,px_495,px_496,px_497,px_498,px_499,px_500,px_501,px_502,px_503,px_504,px_505,px_506,px_507,px_508,px_509,px_510,px_511,px_512,px_513,px_514,px_515,px_516,px_517,px_518,px_519,px_520,px_521,px_522,px_523,px_524,px_525,px_526,px_527,px_528,px_529,px_530,px_531,px_532,px_533,px_534,px_535,px_536,px_537,px_538,px_539,px_540,px_541,px_542,px_543,px_544,px_545,px_546,px_547,px_548,px_549,px_550,px_551,px_552,px_553,px_554,px_555,px_556,px_557,px_558,px_559,px_560,px_561,px_562,px_563,px_564,px_565,px_566,px_567,px_568,px_569,px_570,px_571,px_572,px_573,px_574,px_575,px_576,px_577,px_578,px_579,px_580,px_581,px_582,px_583,px_584,px_585,px_586,px_587,px_588,px_589,px_590,px_591,px_592,px_593,px_594,px_595,px_596,px_597,px_598,px_599,px_600,px_601,px_602,px_603,px_604,px_605,px_606,px_607,px_608,px_609,px_610,px_611,px_612,px_613,px_614,px_615,px_616,px_617,px_618,px_619,px_620,px_621,px_622,px_623,px_624,px_625,px_626,px_627,px_628,px_629,px_630,px_631,px_632,px_633,px_634,px_635,px_636,px_637,px_638,px_639,px_640,px_641,px_642,px_643,px_644,px_645,px_646,px_647,px_648,px_649,px_650,px_651,px_652,px_653,px_654,px_655,px_656,px_657,px_658,px_659,px_660,px_661,px_662,px_663,px_664,px_665,px_666,px_667,px_668,px_669,px_670,px_671,px_672,px_673,px_674,px_675,px_676,px_677,px_678,px_679,px_680,px_681,px_682,px_683,px_684,px_685,px_686,px_687,px_688,px_689,px_690,px_691,px_692,px_693,px_694,px_695,px_696,px_697,px_698,px_699,px_700,px_701,px_702,px_703,px_704,px_705,px_706,px_707,px_708,px_709,px_710,px_711,px_712,px_713,px_714,px_715,px_716,px_717,px_718,px_719,px_720,px_721,px_722,px_723,px_724,px_725,px_726,px_727,px_728,px_729,px_730,px_731,px_732,px_733,px_734,px_735,px_736,px_737,px_738,px_739,px_740,px_741,px_742,px_743,px_744,px_745,px_746,px_747,px_748,px_749,px_750,px_751,px_752,px_753,px_754,px_755,px_756,px_757,px_758,px_759,px_760,px_761,px_762,px_763,px_764,px_765,px_766,px_767,px_768,px_769,px_770,px_771,px_772,px_773,px_774,px_775,px_776,px_777,px_778,px_779,px_780,px_781,px_782,px_783,px_784;

// The possibilies of each number (the final number)
reg [25:0] out_total_0;	// 0
reg [25:0] out_total_1;	// 1
reg [25:0] out_total_2;	// 2
reg [25:0] out_total_3;	// 3
reg [25:0] out_total_4;	// 4
reg [25:0] out_total_5;	// 5
reg [25:0] out_total_6;	// 6
reg [25:0] out_total_7;	// 7
reg [25:0] out_total_8;	// 8
reg [25:0] out_total_9;	// 9	

// The following is the buffer for the multiplier 
wire [9:0] p_0,p_1,p_2,p_3,p_4,p_5,p_6,p_7,p_8,p_9,	p_10,p_11,
           p_12,p_13,p_14,p_15,p_16,p_17,p_18,p_19, p_20,p_21,
		   p_22,p_23,p_24,p_25,p_26,p_27,p_28,p_29, p_30,p_31,
		   p_32,p_33,p_34,p_35,p_36,p_37,p_38,p_39, p_40,p_41,
		   p_42,p_43,p_44,p_45,p_46,p_47,p_48,p_49, p_50,p_51,
		   p_52,p_53,p_54,p_55;
wire [18:0] w_0,w_1,w_2,w_3,w_4,w_5,w_6,w_7,w_8,w_9, w_10,w_11,
            w_12,w_13,w_14,w_15,w_16,w_17,w_18,w_19, w_20,w_21,
			w_22,w_23,w_24,w_25,w_26,w_27,w_28,w_29, w_30,w_31,
			w_32,w_33,w_34,w_35,w_36,w_37,w_38,w_39, w_40,w_41,
			w_42,w_43,w_44,w_45,w_46,w_47,w_48,w_49, w_50,w_51,
			w_52,w_53,w_54,w_55;
reg [9:0] r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,
          r16,r17,r18,r19,r20,r21,r22,r23,r24,r25,r26,r27,r28,r29,
	      r30,r31,r32,r33,r34,r35,r36,r37,r38,r39,r40,r41,r42,r43,
	      r44,r45,r46,r47,r48,r49,r50,r51,r52,r53,r54,r55;
reg [18:0] wr0,wr1,wr2,wr3,wr4,wr5,wr6,wr7,wr8,wr9,wr10,wr11,wr12,
           wr13,wr14,wr15,wr16,wr17,wr18,wr19,wr20,wr21,wr22,wr23,
		   wr24,wr25,wr26,wr27,wr28,wr29,wr30,wr31,wr32,wr33,wr34,
		   wr35,wr36,wr37,wr38,wr39,wr40,wr41,wr42,wr43,wr44,wr45,
		   wr46,wr47,wr48,wr49,wr50,wr51,wr52,wr53,wr54,wr55;

// The following is the buffers for the adder layers
// First layer
wire [25:0] out_temp_0, out_temp_1,out_temp_2,out_temp_3,out_temp_4,out_temp_5,out_temp_6,out_temp_7,out_temp_8,out_temp_9,
		    out_temp_10,out_temp_11,out_temp_12,out_temp_13,out_temp_14,out_temp_15,out_temp_16,out_temp_17,out_temp_18,
			out_temp_19,out_temp_20,out_temp_21,out_temp_22,out_temp_23,out_temp_24,out_temp_25,out_temp_26,out_temp_27,
			out_temp_28,out_temp_29,out_temp_30,out_temp_31,out_temp_32,out_temp_33,out_temp_34,out_temp_35,out_temp_36,
			out_temp_37,out_temp_38,out_temp_39,out_temp_40,out_temp_41,out_temp_42,out_temp_43,out_temp_44,out_temp_45,
			out_temp_46,out_temp_47,out_temp_48,out_temp_49,out_temp_50,out_temp_51,out_temp_52,out_temp_53,out_temp_54,
			out_temp_55;
// Seconde layer
wire [25:0] out_2nd_temp_0,out_2nd_temp_1,out_2nd_temp_2,out_2nd_temp_3,out_2nd_temp_4,out_2nd_temp_5,out_2nd_temp_6,out_2nd_temp_7,
			out_2nd_temp_8,out_2nd_temp_9, out_2nd_temp_10,out_2nd_temp_11,out_2nd_temp_12,out_2nd_temp_13,out_2nd_temp_14,out_2nd_temp_15,
			out_2nd_temp_16,out_2nd_temp_17,out_2nd_temp_18,out_2nd_temp_19, out_2nd_temp_20,out_2nd_temp_21,out_2nd_temp_22,out_2nd_temp_23,
			out_2nd_temp_24,out_2nd_temp_25,out_2nd_temp_26,out_2nd_temp_27; 
// Third layer
wire [25:0] out_3rd_temp_0,out_3rd_temp_1,out_3rd_temp_2,out_3rd_temp_3,out_3rd_temp_4,out_3rd_temp_5,out_3rd_temp_6,out_3rd_temp_7,out_3rd_temp_8,
			out_3rd_temp_9, out_3rd_temp_10,out_3rd_temp_11,out_3rd_temp_12,out_3rd_temp_13;
// Fourth layer
wire [25:0] out_4th_temp_0,out_4th_temp_1,out_4th_temp_2,out_4th_temp_3,out_4th_temp_4,out_4th_temp_5,out_4th_temp_6;
// Fifth layer
wire [25:0] out_5th_temp_0,out_5th_temp_1,out_5th_temp_2,out_5th_temp_3;
// Sixth layer
wire [25:0] out_6th_temp_0,out_6th_temp_1;
// Seventh layer
wire [25:0] out_7th_temp;

// Used to store each output sequence
wire [25:0] out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13;
wire [25:0] temp1,temp2,temp3,temp4,temp5,temp6,temp7,temp_demi;
wire [25:0] temp_2nd_1,temp_2nd_2,temp_2nd_3,temp_2nd_4;
wire [25:0] temp_3rd_1,temp_3rd_2,temp_total,temp_bias;
wire [25:0] temp_output;
//bias wire
wire [18:0] bias_weight;
wire [9:0] bias_pixel;
//register
reg [18:0] bias_w;
reg [9:0] bias_p;
// Buffers for each sequence (784/56)
reg [25:0] out_0; 
reg [25:0] out_1;
reg [25:0] out_2; 
reg [25:0] out_3;
reg [25:0] out_4;
reg [25:0] out_5; 
reg [25:0] out_6;
reg [25:0] out_7;
reg [25:0] out_8; 
reg [25:0] out_9;
reg [25:0] out_10;
reg [25:0] out_11; 
reg [25:0] out_12;
reg [25:0] out_13; 
reg [25:0] out_14;	// Beta

//flag signal
reg [3:0]neuron_flag;

// For case statement
reg [7:0] select;
reg [5:0] state;
reg [4:0] status;
//reg [7:0] seq;
//output_valid
reg ov;
//counter
//reg [5:0] counter;
//reg [3:0] sum_cnt;
//bais wire assignment
assign bias_weight=bias_w;
assign bias_pixel=bias_p;

// Reverse Reset
wire GlobalResetR = ~GlobalReset;
//first iteration flag
reg flag_1st;
//end flag
reg flag_stop;
reg flag_s; //synthsis purpose signal
//reset signal;
reg reset;
reg flagging_neuron;
reg buff;
//mux buffer
reg [25: 0] buffer0;
reg [25: 0] buffer1;
reg [25: 0] buffer2;
reg [25: 0] buffer3;
reg [25: 0] buffer4;
reg [25: 0] buffer5;
reg [25: 0] buffer6;
reg [25: 0] buffer7;
reg [25: 0] buffer8;
reg [25: 0] buffer9;
reg [25: 0] temp_buffer0,temp_buffer1,temp_buffer2,temp_buffer3,temp_buffer4,temp_buffer5,temp_buffer6,temp_buffer7;
reg [25: 0] buffer_select;
reg [3:0] outBuffer;
//output_valid assign
assign Output_Valid=ov;
assign Image_Number=outBuffer;
// Get the value from each input (weight)
assign temp_demi={(25){1'b0}};
assign w_0=wr0;
assign w_1=wr1;
assign w_2=wr2;
assign w_3=wr3;
assign w_4=wr4;
assign w_5=wr5;
assign w_6=wr6;
assign w_7=wr7;
assign w_8=wr8;
assign w_9=wr9;
assign w_10=wr10;
assign w_11=wr11;
assign w_12=wr12;
assign w_13=wr13;
assign w_14=wr14;
assign w_15=wr15;
assign w_16=wr16;
assign w_17=wr17;
assign w_18=wr18;
assign w_19=wr19;
assign w_20=wr20;
assign w_21=wr21;
assign w_22=wr22;
assign w_23=wr23;
assign w_24=wr24;
assign w_25=wr25;
assign w_26=wr26;
assign w_27=wr27;
assign w_28=wr28;
assign w_29=wr29;
assign w_30=wr30;
assign w_31=wr31;
assign w_32=wr32;
assign w_33=wr33;
assign w_34=wr34;
assign w_35=wr35;
assign w_36=wr36;
assign w_37=wr37;
assign w_38=wr38;
assign w_39=wr39;
assign w_40=wr40;
assign w_41=wr41;
assign w_42=wr42;
assign w_43=wr43;
assign w_44=wr44;
assign w_45=wr45;
assign w_46=wr46;
assign w_47=wr47;
assign w_48=wr48;
assign w_49=wr49;
assign w_50=wr50;
assign w_51=wr51;
assign w_52=wr52;
assign w_53=wr53;
assign w_54=wr54;
assign w_55=wr55;

// Get the value from each input (pixel)
assign p_0=r0;
assign p_1=r1;
assign p_2=r2;
assign p_3=r3;
assign p_4=r4;
assign p_5=r5;
assign p_6=r6;
assign p_7=r7;
assign p_8=r8;
assign p_9=r9;
assign p_10=r10;
assign p_11=r11;
assign p_12=r12;
assign p_13=r13;
assign p_14=r14;
assign p_15=r15;
assign p_16=r16;
assign p_17=r17;
assign p_18=r18;
assign p_19=r19;
assign p_20=r20;
assign p_21=r21;
assign p_22=r22;
assign p_23=r23;
assign p_24=r24;
assign p_25=r25;
assign p_26=r26;
assign p_27=r27;
assign p_28=r28;
assign p_29=r29;
assign p_30=r30;
assign p_31=r31;
assign p_32=r32;
assign p_33=r33;
assign p_34=r34;
assign p_35=r35;
assign p_36=r36;
assign p_37=r37;
assign p_38=r38;
assign p_39=r39;
assign p_40=r40;
assign p_41=r41;
assign p_42=r42;
assign p_43=r43;
assign p_44=r44;
assign p_45=r45;
assign p_46=r46;
assign p_47=r47;
assign p_48=r48;
assign p_49=r49;
assign p_50=r50;
assign p_51=r51;
assign p_52=r52;
assign p_53=r53;
assign p_54=r54;
assign p_55=r55;

// Get the result from each sequence
assign out0=out_0;
assign out1=out_1;
assign out2=out_2;
assign out3=out_3;
assign out4=out_4;
assign out5=out_5;
assign out6=out_6;
assign out7=out_7;
assign out8=out_8;
assign out9=out_9;
assign out10=out_10;
assign out11=out_11;
assign out12=out_12;
assign out13=out_13;


// Using 28*2 56 multiplier will do 14 iteration for each neuron
// One more beta add to the summation after each neuron has been calculated
FixedPointMultiplier Multi0(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_0),.PixelPort(p_0),.Output_syn(out_temp_0));//0
FixedPointMultiplier Multi1(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_1),.PixelPort(p_1),.Output_syn(out_temp_1));//1
FixedPointMultiplier Multi2(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_2),.PixelPort(p_2),.Output_syn(out_temp_2));//2
FixedPointMultiplier Multi3(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_3),.PixelPort(p_3),.Output_syn(out_temp_3));//3
FixedPointMultiplier Multi4(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_4),.PixelPort(p_4),.Output_syn(out_temp_4));//4
FixedPointMultiplier Multi5(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_5),.PixelPort(p_5),.Output_syn(out_temp_5));//5
FixedPointMultiplier Multi6(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_6),.PixelPort(p_6),.Output_syn(out_temp_6));//6
FixedPointMultiplier Multi7(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_7),.PixelPort(p_7),.Output_syn(out_temp_7));//7
FixedPointMultiplier Multi8(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_8),.PixelPort(p_8),.Output_syn(out_temp_8));//8
FixedPointMultiplier Multi9(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_9),.PixelPort(p_9),.Output_syn(out_temp_9));//9
FixedPointMultiplier Multi10(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_10),.PixelPort(p_10),.Output_syn(out_temp_10));//10
FixedPointMultiplier Multi11(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_11),.PixelPort(p_11),.Output_syn(out_temp_11));//11
FixedPointMultiplier Multi12(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_12),.PixelPort(p_12),.Output_syn(out_temp_12));//12
FixedPointMultiplier Multi13(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_13),.PixelPort(p_13),.Output_syn(out_temp_13));//13
FixedPointMultiplier Multi14(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_14),.PixelPort(p_14),.Output_syn(out_temp_14));//14
FixedPointMultiplier Multi15(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_15),.PixelPort(p_15),.Output_syn(out_temp_15));//15
FixedPointMultiplier Multi16(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_16),.PixelPort(p_16),.Output_syn(out_temp_16));//16
FixedPointMultiplier Multi17(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_17),.PixelPort(p_17),.Output_syn(out_temp_17));//17
FixedPointMultiplier Multi18(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_18),.PixelPort(p_18),.Output_syn(out_temp_18));//18
FixedPointMultiplier Multi19(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_19),.PixelPort(p_19),.Output_syn(out_temp_19));//19
FixedPointMultiplier Multi20(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_20),.PixelPort(p_20),.Output_syn(out_temp_20));//20
FixedPointMultiplier Multi21(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_21),.PixelPort(p_21),.Output_syn(out_temp_21));//21
FixedPointMultiplier Multi22(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_22),.PixelPort(p_22),.Output_syn(out_temp_22));//22
FixedPointMultiplier Multi23(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_23),.PixelPort(p_23),.Output_syn(out_temp_23));//23
FixedPointMultiplier Multi24(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_24),.PixelPort(p_24),.Output_syn(out_temp_24));//24
FixedPointMultiplier Multi25(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_25),.PixelPort(p_25),.Output_syn(out_temp_25));//25
FixedPointMultiplier Multi26(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_26),.PixelPort(p_26),.Output_syn(out_temp_26));//26
FixedPointMultiplier Multi27(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_27),.PixelPort(p_27),.Output_syn(out_temp_27));//27
FixedPointMultiplier Multi28(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_28),.PixelPort(p_28),.Output_syn(out_temp_28));//28
FixedPointMultiplier Multi29(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_29),.PixelPort(p_29),.Output_syn(out_temp_29));//29
FixedPointMultiplier Multi30(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_30),.PixelPort(p_30),.Output_syn(out_temp_30));//30
FixedPointMultiplier Multi31(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_31),.PixelPort(p_31),.Output_syn(out_temp_31));//31
FixedPointMultiplier Multi32(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_32),.PixelPort(p_32),.Output_syn(out_temp_32));//32
FixedPointMultiplier Multi33(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_33),.PixelPort(p_33),.Output_syn(out_temp_33));//33
FixedPointMultiplier Multi34(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_34),.PixelPort(p_34),.Output_syn(out_temp_34));//34
FixedPointMultiplier Multi35(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_35),.PixelPort(p_35),.Output_syn(out_temp_35));//35
FixedPointMultiplier Multi36(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_36),.PixelPort(p_36),.Output_syn(out_temp_36));//36
FixedPointMultiplier Multi37(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_37),.PixelPort(p_37),.Output_syn(out_temp_37));//37
FixedPointMultiplier Multi38(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_38),.PixelPort(p_38),.Output_syn(out_temp_38));//38
FixedPointMultiplier Multi39(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_39),.PixelPort(p_39),.Output_syn(out_temp_39));//39
FixedPointMultiplier Multi40(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_40),.PixelPort(p_40),.Output_syn(out_temp_40));//40
FixedPointMultiplier Multi41(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_41),.PixelPort(p_41),.Output_syn(out_temp_41));//41
FixedPointMultiplier Multi42(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_42),.PixelPort(p_42),.Output_syn(out_temp_42));//42
FixedPointMultiplier Multi43(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_43),.PixelPort(p_43),.Output_syn(out_temp_43));//43
FixedPointMultiplier Multi44(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_44),.PixelPort(p_44),.Output_syn(out_temp_44));//44
FixedPointMultiplier Multi45(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_45),.PixelPort(p_45),.Output_syn(out_temp_45));//45
FixedPointMultiplier Multi46(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_46),.PixelPort(p_46),.Output_syn(out_temp_46));//46
FixedPointMultiplier Multi47(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_47),.PixelPort(p_47),.Output_syn(out_temp_47));//47
FixedPointMultiplier Multi48(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_48),.PixelPort(p_48),.Output_syn(out_temp_48));//48
FixedPointMultiplier Multi49(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_49),.PixelPort(p_49),.Output_syn(out_temp_49));//49
FixedPointMultiplier Multi50(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_50),.PixelPort(p_50),.Output_syn(out_temp_50));//50
FixedPointMultiplier Multi51(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_51),.PixelPort(p_51),.Output_syn(out_temp_51));//51
FixedPointMultiplier Multi52(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_52),.PixelPort(p_52),.Output_syn(out_temp_52));//52
FixedPointMultiplier Multi53(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_53),.PixelPort(p_53),.Output_syn(out_temp_53));//53
FixedPointMultiplier Multi54(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_54),.PixelPort(p_54),.Output_syn(out_temp_54));//54
FixedPointMultiplier Multi55(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(w_55),.PixelPort(p_55),.Output_syn(out_temp_55));//55

// First layer of adder

FixedPointAdder Addition1_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_0),.Port1(out_temp_1),.Output_syn(out_2nd_temp_0)); //0
FixedPointAdder Addition1_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_2),.Port1(out_temp_3),.Output_syn(out_2nd_temp_1));
FixedPointAdder Addition1_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_4),.Port1(out_temp_5),.Output_syn(out_2nd_temp_2)); //0
FixedPointAdder Addition1_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_6),.Port1(out_temp_7),.Output_syn(out_2nd_temp_3));
FixedPointAdder Addition1_5(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_8),.Port1(out_temp_9),.Output_syn(out_2nd_temp_4)); //0
FixedPointAdder Addition1_6(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_10),.Port1(out_temp_11),.Output_syn(out_2nd_temp_5));
FixedPointAdder Addition1_7(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_12),.Port1(out_temp_13),.Output_syn(out_2nd_temp_6)); //0
FixedPointAdder Addition1_8(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_14),.Port1(out_temp_15),.Output_syn(out_2nd_temp_7));
FixedPointAdder Addition1_9(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_16),.Port1(out_temp_17),.Output_syn(out_2nd_temp_8)); //0
FixedPointAdder Addition1_10(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_18),.Port1(out_temp_19),.Output_syn(out_2nd_temp_9));
FixedPointAdder Addition1_11(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_20),.Port1(out_temp_21),.Output_syn(out_2nd_temp_10)); //0
FixedPointAdder Addition1_12(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_22),.Port1(out_temp_23),.Output_syn(out_2nd_temp_11));
FixedPointAdder Addition1_13(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_24),.Port1(out_temp_25),.Output_syn(out_2nd_temp_12)); //0
FixedPointAdder Addition1_14(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_26),.Port1(out_temp_27),.Output_syn(out_2nd_temp_13));
FixedPointAdder Addition1_15(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_28),.Port1(out_temp_29),.Output_syn(out_2nd_temp_14)); //0
FixedPointAdder Addition1_16(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_30),.Port1(out_temp_31),.Output_syn(out_2nd_temp_15));
FixedPointAdder Addition1_17(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_32),.Port1(out_temp_33),.Output_syn(out_2nd_temp_16)); //0
FixedPointAdder Addition1_18(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_34),.Port1(out_temp_35),.Output_syn(out_2nd_temp_17));
FixedPointAdder Addition1_19(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_36),.Port1(out_temp_37),.Output_syn(out_2nd_temp_18)); //0
FixedPointAdder Addition1_20(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_38),.Port1(out_temp_39),.Output_syn(out_2nd_temp_19));
FixedPointAdder Addition1_21(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_40),.Port1(out_temp_41),.Output_syn(out_2nd_temp_20)); //0
FixedPointAdder Addition1_22(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_42),.Port1(out_temp_43),.Output_syn(out_2nd_temp_21));
FixedPointAdder Addition1_23(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_44),.Port1(out_temp_45),.Output_syn(out_2nd_temp_22)); //0
FixedPointAdder Addition1_24(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_46),.Port1(out_temp_47),.Output_syn(out_2nd_temp_23));
FixedPointAdder Addition1_25(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_48),.Port1(out_temp_49),.Output_syn(out_2nd_temp_24)); //0
FixedPointAdder Addition1_26(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_50),.Port1(out_temp_51),.Output_syn(out_2nd_temp_25));
FixedPointAdder Addition1_27(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_52),.Port1(out_temp_53),.Output_syn(out_2nd_temp_26)); //0
FixedPointAdder Addition1_28(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_temp_54),.Port1(out_temp_55),.Output_syn(out_2nd_temp_27));
//second layer of adder
FixedPointAdder Addition2_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_0),.Port1(out_2nd_temp_1),.Output_syn(out_3rd_temp_0)); 
FixedPointAdder Addition2_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_2),.Port1(out_2nd_temp_3),.Output_syn(out_3rd_temp_1)); 
FixedPointAdder Addition2_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_4),.Port1(out_2nd_temp_5),.Output_syn(out_3rd_temp_2)); 
FixedPointAdder Addition2_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_6),.Port1(out_2nd_temp_7),.Output_syn(out_3rd_temp_3)); 
FixedPointAdder Addition2_5(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_8),.Port1(out_2nd_temp_9),.Output_syn(out_3rd_temp_4)); 
FixedPointAdder Addition2_6(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_10),.Port1(out_2nd_temp_11),.Output_syn(out_3rd_temp_5)); 
FixedPointAdder Addition2_7(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_12),.Port1(out_2nd_temp_13),.Output_syn(out_3rd_temp_6)); 
FixedPointAdder Addition2_8(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_14),.Port1(out_2nd_temp_15),.Output_syn(out_3rd_temp_7)); 
FixedPointAdder Addition2_9(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_16),.Port1(out_2nd_temp_17),.Output_syn(out_3rd_temp_8)); 
FixedPointAdder Addition2_10(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_18),.Port1(out_2nd_temp_19),.Output_syn(out_3rd_temp_9)); 
FixedPointAdder Addition2_11(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_20),.Port1(out_2nd_temp_21),.Output_syn(out_3rd_temp_10)); 
FixedPointAdder Addition2_12(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_22),.Port1(out_2nd_temp_23),.Output_syn(out_3rd_temp_11)); 
FixedPointAdder Addition2_13(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_24),.Port1(out_2nd_temp_25),.Output_syn(out_3rd_temp_12)); 
FixedPointAdder Addition2_14(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_2nd_temp_26),.Port1(out_2nd_temp_27),.Output_syn(out_3rd_temp_13)); 
//third layer of adder
FixedPointAdder Addition3_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_0),.Port1(out_3rd_temp_1),.Output_syn(out_4th_temp_0)); 
FixedPointAdder Addition3_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_2),.Port1(out_3rd_temp_3),.Output_syn(out_4th_temp_1)); 
FixedPointAdder Addition3_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_4),.Port1(out_3rd_temp_5),.Output_syn(out_4th_temp_2)); 
FixedPointAdder Addition3_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_6),.Port1(out_3rd_temp_7),.Output_syn(out_4th_temp_3)); 
FixedPointAdder Addition3_5(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_8),.Port1(out_3rd_temp_9),.Output_syn(out_4th_temp_4)); 
FixedPointAdder Addition3_6(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_10),.Port1(out_3rd_temp_11),.Output_syn(out_4th_temp_5)); 
FixedPointAdder Addition3_7(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_3rd_temp_12),.Port1(out_3rd_temp_13),.Output_syn(out_4th_temp_6)); 
//fourth layer of adder
FixedPointAdder Addition4_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_4th_temp_0),.Port1(out_4th_temp_1),.Output_syn(out_5th_temp_0)); 
FixedPointAdder Addition4_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_4th_temp_2),.Port1(out_4th_temp_3),.Output_syn(out_5th_temp_1)); 
FixedPointAdder Addition4_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_4th_temp_4),.Port1(out_4th_temp_5),.Output_syn(out_5th_temp_2)); 
FixedPointAdder Addition4_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_4th_temp_6),.Port1(temp_demi),.Output_syn(out_5th_temp_3)); //add a demi due to 7 input
//fifth layer
FixedPointAdder Addition5_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_5th_temp_0),.Port1(out_5th_temp_1),.Output_syn(out_6th_temp_0)); 
FixedPointAdder Addition5_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_5th_temp_2),.Port1(out_5th_temp_3),.Output_syn(out_6th_temp_1)); 
//final layer
FixedPointAdder Addition6_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out_6th_temp_0),.Port1(out_6th_temp_1),.Output_syn(out_7th_temp));



//finish 56 multiplication and summation
// Add 14 part together, get each  
FixedPointAdder Addition7_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out0),.Port1(out1),.Output_syn(temp1)); 
FixedPointAdder Addition7_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out2),.Port1(out3),.Output_syn(temp2)); 
FixedPointAdder Addition7_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out4),.Port1(out5),.Output_syn(temp3)); 
FixedPointAdder Addition7_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out6),.Port1(out7),.Output_syn(temp4)); 
FixedPointAdder Addition7_5(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out8),.Port1(out9),.Output_syn(temp5)); 
FixedPointAdder Addition7_6(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out10),.Port1(out11),.Output_syn(temp6)); 
FixedPointAdder Addition7_7(.clk(clk),.GlobalReset(GlobalResetR),.Port2(out12),.Port1(out13),.Output_syn(temp7)); 
FixedPointAdder Addition8_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp1),.Port1(temp2),.Output_syn(temp_2nd_1)); 
FixedPointAdder Addition8_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp3),.Port1(temp4),.Output_syn(temp_2nd_2)); 
FixedPointAdder Addition8_3(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp5),.Port1(temp6),.Output_syn(temp_2nd_3)); 
FixedPointAdder Addition8_4(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp7),.Port1(temp_demi),.Output_syn(temp_2nd_4)); 
FixedPointAdder Addition9_1(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp_2nd_1),.Port1(temp_2nd_2),.Output_syn(temp_3rd_1)); 
FixedPointAdder Addition9_2(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp_2nd_3),.Port1(temp_2nd_4),.Output_syn(temp_3rd_2)); 
FixedPointAdder Addition10(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp_3rd_1),.Port1(temp_3rd_2),.Output_syn(temp_total)); 

//bias
FixedPointMultiplier Multibias(.clk(clk),.GlobalReset(GlobalResetR),.WeightPort(bias_weight),.PixelPort(bias_pixel),.Output_syn(temp_bias));//bias
FixedPointAdder Additionb(.clk(clk),.GlobalReset(GlobalResetR),.Port2(temp_total),.Port1(temp_bias),.Output_syn(temp_output)); 

always @(posedge clk or negedge GlobalReset) begin
	if (GlobalReset == 1'b0)
		begin
			//select <= 0;
		end
	else
		begin
			if(Input_Valid)
				begin
					//input all pixel value
					px_0<=Pix_0; px_1<=Pix_1; px_2<=Pix_2; px_3<=Pix_3; px_4<=Pix_4; px_5<=Pix_5; px_6<=Pix_6; px_7<=Pix_7; px_8<=Pix_8; px_9<=Pix_9; px_10<=Pix_10; px_11<=Pix_11; px_12<=Pix_12; px_13<=Pix_13; px_14<=Pix_14; px_15<=Pix_15; px_16<=Pix_16; px_17<=Pix_17; px_18<=Pix_18; px_19<=Pix_19; px_20<=Pix_20; px_21<=Pix_21; px_22<=Pix_22; px_23<=Pix_23; px_24<=Pix_24; px_25<=Pix_25; px_26<=Pix_26; px_27<=Pix_27; px_28<=Pix_28; px_29<=Pix_29; px_30<=Pix_30; px_31<=Pix_31; px_32<=Pix_32; px_33<=Pix_33; px_34<=Pix_34; px_35<=Pix_35; px_36<=Pix_36; px_37<=Pix_37; px_38<=Pix_38; px_39<=Pix_39; px_40<=Pix_40; px_41<=Pix_41; px_42<=Pix_42; px_43<=Pix_43; px_44<=Pix_44; px_45<=Pix_45; px_46<=Pix_46; px_47<=Pix_47; px_48<=Pix_48; px_49<=Pix_49; px_50<=Pix_50; px_51<=Pix_51; px_52<=Pix_52; px_53<=Pix_53; px_54<=Pix_54; px_55<=Pix_55; px_56<=Pix_56; px_57<=Pix_57; px_58<=Pix_58; px_59<=Pix_59; px_60<=Pix_60; px_61<=Pix_61; px_62<=Pix_62; px_63<=Pix_63; px_64<=Pix_64; px_65<=Pix_65; px_66<=Pix_66; px_67<=Pix_67; px_68<=Pix_68; px_69<=Pix_69; px_70<=Pix_70; px_71<=Pix_71; px_72<=Pix_72; px_73<=Pix_73; px_74<=Pix_74; px_75<=Pix_75; px_76<=Pix_76; px_77<=Pix_77; px_78<=Pix_78; px_79<=Pix_79; px_80<=Pix_80; px_81<=Pix_81; px_82<=Pix_82; px_83<=Pix_83; px_84<=Pix_84; px_85<=Pix_85; px_86<=Pix_86; px_87<=Pix_87; px_88<=Pix_88; px_89<=Pix_89; px_90<=Pix_90; px_91<=Pix_91; px_92<=Pix_92; px_93<=Pix_93; px_94<=Pix_94; px_95<=Pix_95; px_96<=Pix_96; px_97<=Pix_97; px_98<=Pix_98; px_99<=Pix_99; px_100<=Pix_100; px_101<=Pix_101; px_102<=Pix_102; px_103<=Pix_103; px_104<=Pix_104; px_105<=Pix_105; px_106<=Pix_106; px_107<=Pix_107; px_108<=Pix_108; px_109<=Pix_109; px_110<=Pix_110; px_111<=Pix_111; px_112<=Pix_112; px_113<=Pix_113; px_114<=Pix_114; px_115<=Pix_115; px_116<=Pix_116; px_117<=Pix_117; px_118<=Pix_118; px_119<=Pix_119; px_120<=Pix_120; px_121<=Pix_121; px_122<=Pix_122; px_123<=Pix_123; px_124<=Pix_124; px_125<=Pix_125; px_126<=Pix_126; px_127<=Pix_127; px_128<=Pix_128; px_129<=Pix_129; px_130<=Pix_130; px_131<=Pix_131; px_132<=Pix_132; px_133<=Pix_133; px_134<=Pix_134; px_135<=Pix_135; px_136<=Pix_136; px_137<=Pix_137; px_138<=Pix_138; px_139<=Pix_139; px_140<=Pix_140; px_141<=Pix_141; px_142<=Pix_142; px_143<=Pix_143; px_144<=Pix_144; px_145<=Pix_145; px_146<=Pix_146; px_147<=Pix_147; px_148<=Pix_148; px_149<=Pix_149; px_150<=Pix_150; px_151<=Pix_151; px_152<=Pix_152; px_153<=Pix_153; px_154<=Pix_154; px_155<=Pix_155; px_156<=Pix_156; px_157<=Pix_157; px_158<=Pix_158; px_159<=Pix_159; px_160<=Pix_160; px_161<=Pix_161; px_162<=Pix_162; px_163<=Pix_163; px_164<=Pix_164; px_165<=Pix_165; px_166<=Pix_166; px_167<=Pix_167; px_168<=Pix_168; px_169<=Pix_169; px_170<=Pix_170; px_171<=Pix_171; px_172<=Pix_172; px_173<=Pix_173; px_174<=Pix_174; px_175<=Pix_175; px_176<=Pix_176; px_177<=Pix_177; px_178<=Pix_178; px_179<=Pix_179; px_180<=Pix_180; px_181<=Pix_181; px_182<=Pix_182; px_183<=Pix_183; px_184<=Pix_184; px_185<=Pix_185; px_186<=Pix_186; px_187<=Pix_187; px_188<=Pix_188; px_189<=Pix_189; px_190<=Pix_190; px_191<=Pix_191; px_192<=Pix_192; px_193<=Pix_193; px_194<=Pix_194; px_195<=Pix_195; px_196<=Pix_196; px_197<=Pix_197; px_198<=Pix_198; px_199<=Pix_199; px_200<=Pix_200; px_201<=Pix_201; px_202<=Pix_202; px_203<=Pix_203; px_204<=Pix_204; px_205<=Pix_205; px_206<=Pix_206; px_207<=Pix_207; px_208<=Pix_208; px_209<=Pix_209; px_210<=Pix_210; px_211<=Pix_211; px_212<=Pix_212; px_213<=Pix_213; px_214<=Pix_214; px_215<=Pix_215; px_216<=Pix_216; px_217<=Pix_217; px_218<=Pix_218; px_219<=Pix_219; px_220<=Pix_220; px_221<=Pix_221; px_222<=Pix_222; px_223<=Pix_223; px_224<=Pix_224; px_225<=Pix_225; px_226<=Pix_226; px_227<=Pix_227; px_228<=Pix_228; px_229<=Pix_229; px_230<=Pix_230; px_231<=Pix_231; px_232<=Pix_232; px_233<=Pix_233; px_234<=Pix_234; px_235<=Pix_235; px_236<=Pix_236; px_237<=Pix_237; px_238<=Pix_238; px_239<=Pix_239; px_240<=Pix_240; px_241<=Pix_241; px_242<=Pix_242; px_243<=Pix_243; px_244<=Pix_244; px_245<=Pix_245; px_246<=Pix_246; px_247<=Pix_247; px_248<=Pix_248; px_249<=Pix_249; px_250<=Pix_250; px_251<=Pix_251; px_252<=Pix_252; px_253<=Pix_253; px_254<=Pix_254; px_255<=Pix_255; px_256<=Pix_256; px_257<=Pix_257; px_258<=Pix_258; px_259<=Pix_259; px_260<=Pix_260; px_261<=Pix_261; px_262<=Pix_262; px_263<=Pix_263; px_264<=Pix_264; px_265<=Pix_265; px_266<=Pix_266; px_267<=Pix_267; px_268<=Pix_268; px_269<=Pix_269; px_270<=Pix_270; px_271<=Pix_271; px_272<=Pix_272; px_273<=Pix_273; px_274<=Pix_274; px_275<=Pix_275; px_276<=Pix_276; px_277<=Pix_277; px_278<=Pix_278; px_279<=Pix_279; px_280<=Pix_280; px_281<=Pix_281; px_282<=Pix_282; px_283<=Pix_283; px_284<=Pix_284; px_285<=Pix_285; px_286<=Pix_286; px_287<=Pix_287; px_288<=Pix_288; px_289<=Pix_289; px_290<=Pix_290; px_291<=Pix_291; px_292<=Pix_292; px_293<=Pix_293; px_294<=Pix_294; px_295<=Pix_295; px_296<=Pix_296; px_297<=Pix_297; px_298<=Pix_298; px_299<=Pix_299; px_300<=Pix_300; px_301<=Pix_301; px_302<=Pix_302; px_303<=Pix_303; px_304<=Pix_304; px_305<=Pix_305; px_306<=Pix_306; px_307<=Pix_307; px_308<=Pix_308; px_309<=Pix_309; px_310<=Pix_310; px_311<=Pix_311; px_312<=Pix_312; px_313<=Pix_313; px_314<=Pix_314; px_315<=Pix_315; px_316<=Pix_316; px_317<=Pix_317; px_318<=Pix_318; px_319<=Pix_319; px_320<=Pix_320; px_321<=Pix_321; px_322<=Pix_322; px_323<=Pix_323; px_324<=Pix_324; px_325<=Pix_325; px_326<=Pix_326; px_327<=Pix_327; px_328<=Pix_328; px_329<=Pix_329; px_330<=Pix_330; px_331<=Pix_331; px_332<=Pix_332; px_333<=Pix_333; px_334<=Pix_334; px_335<=Pix_335; px_336<=Pix_336; px_337<=Pix_337; px_338<=Pix_338; px_339<=Pix_339; px_340<=Pix_340; px_341<=Pix_341; px_342<=Pix_342; px_343<=Pix_343; px_344<=Pix_344; px_345<=Pix_345; px_346<=Pix_346; px_347<=Pix_347; px_348<=Pix_348; px_349<=Pix_349; px_350<=Pix_350; px_351<=Pix_351; px_352<=Pix_352; px_353<=Pix_353; px_354<=Pix_354; px_355<=Pix_355; px_356<=Pix_356; px_357<=Pix_357; px_358<=Pix_358; px_359<=Pix_359; px_360<=Pix_360; px_361<=Pix_361; px_362<=Pix_362; px_363<=Pix_363; px_364<=Pix_364; px_365<=Pix_365; px_366<=Pix_366; px_367<=Pix_367; px_368<=Pix_368; px_369<=Pix_369; px_370<=Pix_370; px_371<=Pix_371; px_372<=Pix_372; px_373<=Pix_373; px_374<=Pix_374; px_375<=Pix_375; px_376<=Pix_376; px_377<=Pix_377; px_378<=Pix_378; px_379<=Pix_379; px_380<=Pix_380; px_381<=Pix_381; px_382<=Pix_382; px_383<=Pix_383; px_384<=Pix_384; px_385<=Pix_385; px_386<=Pix_386; px_387<=Pix_387; px_388<=Pix_388; px_389<=Pix_389; px_390<=Pix_390; px_391<=Pix_391; px_392<=Pix_392; px_393<=Pix_393; px_394<=Pix_394; px_395<=Pix_395; px_396<=Pix_396; px_397<=Pix_397; px_398<=Pix_398; px_399<=Pix_399; px_400<=Pix_400; px_401<=Pix_401; px_402<=Pix_402; px_403<=Pix_403; px_404<=Pix_404; px_405<=Pix_405; px_406<=Pix_406; px_407<=Pix_407; px_408<=Pix_408; px_409<=Pix_409; px_410<=Pix_410; px_411<=Pix_411; px_412<=Pix_412; px_413<=Pix_413; px_414<=Pix_414; px_415<=Pix_415; px_416<=Pix_416; px_417<=Pix_417; px_418<=Pix_418; px_419<=Pix_419; px_420<=Pix_420; px_421<=Pix_421; px_422<=Pix_422; px_423<=Pix_423; px_424<=Pix_424; px_425<=Pix_425; px_426<=Pix_426; px_427<=Pix_427; px_428<=Pix_428; px_429<=Pix_429; px_430<=Pix_430; px_431<=Pix_431; px_432<=Pix_432; px_433<=Pix_433; px_434<=Pix_434; px_435<=Pix_435; px_436<=Pix_436; px_437<=Pix_437; px_438<=Pix_438; px_439<=Pix_439; px_440<=Pix_440; px_441<=Pix_441; px_442<=Pix_442; px_443<=Pix_443; px_444<=Pix_444; px_445<=Pix_445; px_446<=Pix_446; px_447<=Pix_447; px_448<=Pix_448; px_449<=Pix_449; px_450<=Pix_450; px_451<=Pix_451; px_452<=Pix_452; px_453<=Pix_453; px_454<=Pix_454; px_455<=Pix_455; px_456<=Pix_456; px_457<=Pix_457; px_458<=Pix_458; px_459<=Pix_459; px_460<=Pix_460; px_461<=Pix_461; px_462<=Pix_462; px_463<=Pix_463; px_464<=Pix_464; px_465<=Pix_465; px_466<=Pix_466; px_467<=Pix_467; px_468<=Pix_468; px_469<=Pix_469; px_470<=Pix_470; px_471<=Pix_471; px_472<=Pix_472; px_473<=Pix_473; px_474<=Pix_474; px_475<=Pix_475; px_476<=Pix_476; px_477<=Pix_477; px_478<=Pix_478; px_479<=Pix_479; px_480<=Pix_480; px_481<=Pix_481; px_482<=Pix_482; px_483<=Pix_483; px_484<=Pix_484; px_485<=Pix_485; px_486<=Pix_486; px_487<=Pix_487; px_488<=Pix_488; px_489<=Pix_489; px_490<=Pix_490; px_491<=Pix_491; px_492<=Pix_492; px_493<=Pix_493; px_494<=Pix_494; px_495<=Pix_495; px_496<=Pix_496; px_497<=Pix_497; px_498<=Pix_498; px_499<=Pix_499; px_500<=Pix_500; px_501<=Pix_501; px_502<=Pix_502; px_503<=Pix_503; px_504<=Pix_504; px_505<=Pix_505; px_506<=Pix_506; px_507<=Pix_507; px_508<=Pix_508; px_509<=Pix_509; px_510<=Pix_510; px_511<=Pix_511; px_512<=Pix_512; px_513<=Pix_513; px_514<=Pix_514; px_515<=Pix_515; px_516<=Pix_516; px_517<=Pix_517; px_518<=Pix_518; px_519<=Pix_519; px_520<=Pix_520; px_521<=Pix_521; px_522<=Pix_522; px_523<=Pix_523; px_524<=Pix_524; px_525<=Pix_525; px_526<=Pix_526; px_527<=Pix_527; px_528<=Pix_528; px_529<=Pix_529; px_530<=Pix_530; px_531<=Pix_531; px_532<=Pix_532; px_533<=Pix_533; px_534<=Pix_534; px_535<=Pix_535; px_536<=Pix_536; px_537<=Pix_537; px_538<=Pix_538; px_539<=Pix_539; px_540<=Pix_540; px_541<=Pix_541; px_542<=Pix_542; px_543<=Pix_543; px_544<=Pix_544; px_545<=Pix_545; px_546<=Pix_546; px_547<=Pix_547; px_548<=Pix_548; px_549<=Pix_549; px_550<=Pix_550; px_551<=Pix_551; px_552<=Pix_552; px_553<=Pix_553; px_554<=Pix_554; px_555<=Pix_555; px_556<=Pix_556; px_557<=Pix_557; px_558<=Pix_558; px_559<=Pix_559; px_560<=Pix_560; px_561<=Pix_561; px_562<=Pix_562; px_563<=Pix_563; px_564<=Pix_564; px_565<=Pix_565; px_566<=Pix_566; px_567<=Pix_567; px_568<=Pix_568; px_569<=Pix_569; px_570<=Pix_570; px_571<=Pix_571; px_572<=Pix_572; px_573<=Pix_573; px_574<=Pix_574; px_575<=Pix_575; px_576<=Pix_576; px_577<=Pix_577; px_578<=Pix_578; px_579<=Pix_579; px_580<=Pix_580; px_581<=Pix_581; px_582<=Pix_582; px_583<=Pix_583; px_584<=Pix_584; px_585<=Pix_585; px_586<=Pix_586; px_587<=Pix_587; px_588<=Pix_588; px_589<=Pix_589; px_590<=Pix_590; px_591<=Pix_591; px_592<=Pix_592; px_593<=Pix_593; px_594<=Pix_594; px_595<=Pix_595; px_596<=Pix_596; px_597<=Pix_597; px_598<=Pix_598; px_599<=Pix_599; px_600<=Pix_600; px_601<=Pix_601; px_602<=Pix_602; px_603<=Pix_603; px_604<=Pix_604; px_605<=Pix_605; px_606<=Pix_606; px_607<=Pix_607; px_608<=Pix_608; px_609<=Pix_609; px_610<=Pix_610; px_611<=Pix_611; px_612<=Pix_612; px_613<=Pix_613; px_614<=Pix_614; px_615<=Pix_615; px_616<=Pix_616; px_617<=Pix_617; px_618<=Pix_618; px_619<=Pix_619; px_620<=Pix_620; px_621<=Pix_621; px_622<=Pix_622; px_623<=Pix_623; px_624<=Pix_624; px_625<=Pix_625; px_626<=Pix_626; px_627<=Pix_627; px_628<=Pix_628; px_629<=Pix_629; px_630<=Pix_630; px_631<=Pix_631; px_632<=Pix_632; px_633<=Pix_633; px_634<=Pix_634; px_635<=Pix_635; px_636<=Pix_636; px_637<=Pix_637; px_638<=Pix_638; px_639<=Pix_639; px_640<=Pix_640; px_641<=Pix_641; px_642<=Pix_642; px_643<=Pix_643; px_644<=Pix_644; px_645<=Pix_645; px_646<=Pix_646; px_647<=Pix_647; px_648<=Pix_648; px_649<=Pix_649; px_650<=Pix_650; px_651<=Pix_651; px_652<=Pix_652; px_653<=Pix_653; px_654<=Pix_654; px_655<=Pix_655; px_656<=Pix_656; px_657<=Pix_657; px_658<=Pix_658; px_659<=Pix_659; px_660<=Pix_660; px_661<=Pix_661; px_662<=Pix_662; px_663<=Pix_663; px_664<=Pix_664; px_665<=Pix_665; px_666<=Pix_666; px_667<=Pix_667; px_668<=Pix_668; px_669<=Pix_669; px_670<=Pix_670; px_671<=Pix_671; px_672<=Pix_672; px_673<=Pix_673; px_674<=Pix_674; px_675<=Pix_675; px_676<=Pix_676; px_677<=Pix_677; px_678<=Pix_678; px_679<=Pix_679; px_680<=Pix_680; px_681<=Pix_681; px_682<=Pix_682; px_683<=Pix_683; px_684<=Pix_684; px_685<=Pix_685; px_686<=Pix_686; px_687<=Pix_687; px_688<=Pix_688; px_689<=Pix_689; px_690<=Pix_690; px_691<=Pix_691; px_692<=Pix_692; px_693<=Pix_693; px_694<=Pix_694; px_695<=Pix_695; px_696<=Pix_696; px_697<=Pix_697; px_698<=Pix_698; px_699<=Pix_699; px_700<=Pix_700; px_701<=Pix_701; px_702<=Pix_702; px_703<=Pix_703; px_704<=Pix_704; px_705<=Pix_705; px_706<=Pix_706; px_707<=Pix_707; px_708<=Pix_708; px_709<=Pix_709; px_710<=Pix_710; px_711<=Pix_711; px_712<=Pix_712; px_713<=Pix_713; px_714<=Pix_714; px_715<=Pix_715; px_716<=Pix_716; px_717<=Pix_717; px_718<=Pix_718; px_719<=Pix_719; px_720<=Pix_720; px_721<=Pix_721; px_722<=Pix_722; px_723<=Pix_723; px_724<=Pix_724; px_725<=Pix_725; px_726<=Pix_726; px_727<=Pix_727; px_728<=Pix_728; px_729<=Pix_729; px_730<=Pix_730; px_731<=Pix_731; px_732<=Pix_732; px_733<=Pix_733; px_734<=Pix_734; px_735<=Pix_735; px_736<=Pix_736; px_737<=Pix_737; px_738<=Pix_738; px_739<=Pix_739; px_740<=Pix_740; px_741<=Pix_741; px_742<=Pix_742; px_743<=Pix_743; px_744<=Pix_744; px_745<=Pix_745; px_746<=Pix_746; px_747<=Pix_747; px_748<=Pix_748; px_749<=Pix_749; px_750<=Pix_750; px_751<=Pix_751; px_752<=Pix_752; px_753<=Pix_753; px_754<=Pix_754; px_755<=Pix_755; px_756<=Pix_756; px_757<=Pix_757; px_758<=Pix_758; px_759<=Pix_759; px_760<=Pix_760; px_761<=Pix_761; px_762<=Pix_762; px_763<=Pix_763; px_764<=Pix_764; px_765<=Pix_765; px_766<=Pix_766; px_767<=Pix_767; px_768<=Pix_768; px_769<=Pix_769; px_770<=Pix_770; px_771<=Pix_771; px_772<=Pix_772; px_773<=Pix_773; px_774<=Pix_774; px_775<=Pix_775; px_776<=Pix_776; px_777<=Pix_777; px_778<=Pix_778; px_779<=Pix_779; px_780<=Pix_780; px_781<=Pix_781; px_782<=Pix_782; px_783<=Pix_783; px_784<=Pix_784;  
					w_0_0<=Wgt_0_0; w_0_1<=Wgt_0_1; w_0_2<=Wgt_0_2; w_0_3<=Wgt_0_3; w_0_4<=Wgt_0_4; w_0_5<=Wgt_0_5; w_0_6<=Wgt_0_6; w_0_7<=Wgt_0_7; w_0_8<=Wgt_0_8; w_0_9<=Wgt_0_9; w_0_10<=Wgt_0_10; w_0_11<=Wgt_0_11; w_0_12<=Wgt_0_12; w_0_13<=Wgt_0_13; w_0_14<=Wgt_0_14; w_0_15<=Wgt_0_15; w_0_16<=Wgt_0_16; w_0_17<=Wgt_0_17; w_0_18<=Wgt_0_18; w_0_19<=Wgt_0_19; w_0_20<=Wgt_0_20; w_0_21<=Wgt_0_21; w_0_22<=Wgt_0_22; w_0_23<=Wgt_0_23; w_0_24<=Wgt_0_24; w_0_25<=Wgt_0_25; w_0_26<=Wgt_0_26; w_0_27<=Wgt_0_27; w_0_28<=Wgt_0_28; w_0_29<=Wgt_0_29; w_0_30<=Wgt_0_30; w_0_31<=Wgt_0_31; w_0_32<=Wgt_0_32; w_0_33<=Wgt_0_33; w_0_34<=Wgt_0_34; w_0_35<=Wgt_0_35; w_0_36<=Wgt_0_36; w_0_37<=Wgt_0_37; w_0_38<=Wgt_0_38; w_0_39<=Wgt_0_39; w_0_40<=Wgt_0_40; w_0_41<=Wgt_0_41; w_0_42<=Wgt_0_42; w_0_43<=Wgt_0_43; w_0_44<=Wgt_0_44; w_0_45<=Wgt_0_45; w_0_46<=Wgt_0_46; w_0_47<=Wgt_0_47; w_0_48<=Wgt_0_48; w_0_49<=Wgt_0_49; w_0_50<=Wgt_0_50; w_0_51<=Wgt_0_51; w_0_52<=Wgt_0_52; w_0_53<=Wgt_0_53; w_0_54<=Wgt_0_54; w_0_55<=Wgt_0_55; w_0_56<=Wgt_0_56; w_0_57<=Wgt_0_57; w_0_58<=Wgt_0_58; w_0_59<=Wgt_0_59; w_0_60<=Wgt_0_60; w_0_61<=Wgt_0_61; w_0_62<=Wgt_0_62; w_0_63<=Wgt_0_63; w_0_64<=Wgt_0_64; w_0_65<=Wgt_0_65; w_0_66<=Wgt_0_66; w_0_67<=Wgt_0_67; w_0_68<=Wgt_0_68; w_0_69<=Wgt_0_69; w_0_70<=Wgt_0_70; w_0_71<=Wgt_0_71; w_0_72<=Wgt_0_72; w_0_73<=Wgt_0_73; w_0_74<=Wgt_0_74; w_0_75<=Wgt_0_75; w_0_76<=Wgt_0_76; w_0_77<=Wgt_0_77; w_0_78<=Wgt_0_78; w_0_79<=Wgt_0_79; w_0_80<=Wgt_0_80; w_0_81<=Wgt_0_81; w_0_82<=Wgt_0_82; w_0_83<=Wgt_0_83; w_0_84<=Wgt_0_84; w_0_85<=Wgt_0_85; w_0_86<=Wgt_0_86; w_0_87<=Wgt_0_87; w_0_88<=Wgt_0_88; w_0_89<=Wgt_0_89; w_0_90<=Wgt_0_90; w_0_91<=Wgt_0_91; w_0_92<=Wgt_0_92; w_0_93<=Wgt_0_93; w_0_94<=Wgt_0_94; w_0_95<=Wgt_0_95; w_0_96<=Wgt_0_96; w_0_97<=Wgt_0_97; w_0_98<=Wgt_0_98; w_0_99<=Wgt_0_99; w_0_100<=Wgt_0_100; w_0_101<=Wgt_0_101; w_0_102<=Wgt_0_102; w_0_103<=Wgt_0_103; w_0_104<=Wgt_0_104; w_0_105<=Wgt_0_105; w_0_106<=Wgt_0_106; w_0_107<=Wgt_0_107; w_0_108<=Wgt_0_108; w_0_109<=Wgt_0_109; w_0_110<=Wgt_0_110; w_0_111<=Wgt_0_111; w_0_112<=Wgt_0_112; w_0_113<=Wgt_0_113; w_0_114<=Wgt_0_114; w_0_115<=Wgt_0_115; w_0_116<=Wgt_0_116; w_0_117<=Wgt_0_117; w_0_118<=Wgt_0_118; w_0_119<=Wgt_0_119; w_0_120<=Wgt_0_120; w_0_121<=Wgt_0_121; w_0_122<=Wgt_0_122; w_0_123<=Wgt_0_123; w_0_124<=Wgt_0_124; w_0_125<=Wgt_0_125; w_0_126<=Wgt_0_126; w_0_127<=Wgt_0_127; w_0_128<=Wgt_0_128; w_0_129<=Wgt_0_129; w_0_130<=Wgt_0_130; w_0_131<=Wgt_0_131; w_0_132<=Wgt_0_132; w_0_133<=Wgt_0_133; w_0_134<=Wgt_0_134; w_0_135<=Wgt_0_135; w_0_136<=Wgt_0_136; w_0_137<=Wgt_0_137; w_0_138<=Wgt_0_138; w_0_139<=Wgt_0_139; w_0_140<=Wgt_0_140; w_0_141<=Wgt_0_141; w_0_142<=Wgt_0_142; w_0_143<=Wgt_0_143; w_0_144<=Wgt_0_144; w_0_145<=Wgt_0_145; w_0_146<=Wgt_0_146; w_0_147<=Wgt_0_147; w_0_148<=Wgt_0_148; w_0_149<=Wgt_0_149; w_0_150<=Wgt_0_150; w_0_151<=Wgt_0_151; w_0_152<=Wgt_0_152; w_0_153<=Wgt_0_153; w_0_154<=Wgt_0_154; w_0_155<=Wgt_0_155; w_0_156<=Wgt_0_156; w_0_157<=Wgt_0_157; w_0_158<=Wgt_0_158; w_0_159<=Wgt_0_159; w_0_160<=Wgt_0_160; w_0_161<=Wgt_0_161; w_0_162<=Wgt_0_162; w_0_163<=Wgt_0_163; w_0_164<=Wgt_0_164; w_0_165<=Wgt_0_165; w_0_166<=Wgt_0_166; w_0_167<=Wgt_0_167; w_0_168<=Wgt_0_168; w_0_169<=Wgt_0_169; w_0_170<=Wgt_0_170; w_0_171<=Wgt_0_171; w_0_172<=Wgt_0_172; w_0_173<=Wgt_0_173; w_0_174<=Wgt_0_174; w_0_175<=Wgt_0_175; w_0_176<=Wgt_0_176; w_0_177<=Wgt_0_177; w_0_178<=Wgt_0_178; w_0_179<=Wgt_0_179; w_0_180<=Wgt_0_180; w_0_181<=Wgt_0_181; w_0_182<=Wgt_0_182; w_0_183<=Wgt_0_183; w_0_184<=Wgt_0_184; w_0_185<=Wgt_0_185; w_0_186<=Wgt_0_186; w_0_187<=Wgt_0_187; w_0_188<=Wgt_0_188; w_0_189<=Wgt_0_189; w_0_190<=Wgt_0_190; w_0_191<=Wgt_0_191; w_0_192<=Wgt_0_192; w_0_193<=Wgt_0_193; w_0_194<=Wgt_0_194; w_0_195<=Wgt_0_195; w_0_196<=Wgt_0_196; w_0_197<=Wgt_0_197; w_0_198<=Wgt_0_198; w_0_199<=Wgt_0_199; w_0_200<=Wgt_0_200; w_0_201<=Wgt_0_201; w_0_202<=Wgt_0_202; w_0_203<=Wgt_0_203; w_0_204<=Wgt_0_204; w_0_205<=Wgt_0_205; w_0_206<=Wgt_0_206; w_0_207<=Wgt_0_207; w_0_208<=Wgt_0_208; w_0_209<=Wgt_0_209; w_0_210<=Wgt_0_210; w_0_211<=Wgt_0_211; w_0_212<=Wgt_0_212; w_0_213<=Wgt_0_213; w_0_214<=Wgt_0_214; w_0_215<=Wgt_0_215; w_0_216<=Wgt_0_216; w_0_217<=Wgt_0_217; w_0_218<=Wgt_0_218; w_0_219<=Wgt_0_219; w_0_220<=Wgt_0_220; w_0_221<=Wgt_0_221; w_0_222<=Wgt_0_222; w_0_223<=Wgt_0_223; w_0_224<=Wgt_0_224; w_0_225<=Wgt_0_225; w_0_226<=Wgt_0_226; w_0_227<=Wgt_0_227; w_0_228<=Wgt_0_228; w_0_229<=Wgt_0_229; w_0_230<=Wgt_0_230; w_0_231<=Wgt_0_231; w_0_232<=Wgt_0_232; w_0_233<=Wgt_0_233; w_0_234<=Wgt_0_234; w_0_235<=Wgt_0_235; w_0_236<=Wgt_0_236; w_0_237<=Wgt_0_237; w_0_238<=Wgt_0_238; w_0_239<=Wgt_0_239; w_0_240<=Wgt_0_240; w_0_241<=Wgt_0_241; w_0_242<=Wgt_0_242; w_0_243<=Wgt_0_243; w_0_244<=Wgt_0_244; w_0_245<=Wgt_0_245; w_0_246<=Wgt_0_246; w_0_247<=Wgt_0_247; w_0_248<=Wgt_0_248; w_0_249<=Wgt_0_249; w_0_250<=Wgt_0_250; w_0_251<=Wgt_0_251; w_0_252<=Wgt_0_252; w_0_253<=Wgt_0_253; w_0_254<=Wgt_0_254; w_0_255<=Wgt_0_255; w_0_256<=Wgt_0_256; w_0_257<=Wgt_0_257; w_0_258<=Wgt_0_258; w_0_259<=Wgt_0_259; w_0_260<=Wgt_0_260; w_0_261<=Wgt_0_261; w_0_262<=Wgt_0_262; w_0_263<=Wgt_0_263; w_0_264<=Wgt_0_264; w_0_265<=Wgt_0_265; w_0_266<=Wgt_0_266; w_0_267<=Wgt_0_267; w_0_268<=Wgt_0_268; w_0_269<=Wgt_0_269; w_0_270<=Wgt_0_270; w_0_271<=Wgt_0_271; w_0_272<=Wgt_0_272; w_0_273<=Wgt_0_273; w_0_274<=Wgt_0_274; w_0_275<=Wgt_0_275; w_0_276<=Wgt_0_276; w_0_277<=Wgt_0_277; w_0_278<=Wgt_0_278; w_0_279<=Wgt_0_279; w_0_280<=Wgt_0_280; w_0_281<=Wgt_0_281; w_0_282<=Wgt_0_282; w_0_283<=Wgt_0_283; w_0_284<=Wgt_0_284; w_0_285<=Wgt_0_285; w_0_286<=Wgt_0_286; w_0_287<=Wgt_0_287; w_0_288<=Wgt_0_288; w_0_289<=Wgt_0_289; w_0_290<=Wgt_0_290; w_0_291<=Wgt_0_291; w_0_292<=Wgt_0_292; w_0_293<=Wgt_0_293; w_0_294<=Wgt_0_294; w_0_295<=Wgt_0_295; w_0_296<=Wgt_0_296; w_0_297<=Wgt_0_297; w_0_298<=Wgt_0_298; w_0_299<=Wgt_0_299; w_0_300<=Wgt_0_300; w_0_301<=Wgt_0_301; w_0_302<=Wgt_0_302; w_0_303<=Wgt_0_303; w_0_304<=Wgt_0_304; w_0_305<=Wgt_0_305; w_0_306<=Wgt_0_306; w_0_307<=Wgt_0_307; w_0_308<=Wgt_0_308; w_0_309<=Wgt_0_309; w_0_310<=Wgt_0_310; w_0_311<=Wgt_0_311; w_0_312<=Wgt_0_312; w_0_313<=Wgt_0_313; w_0_314<=Wgt_0_314; w_0_315<=Wgt_0_315; w_0_316<=Wgt_0_316; w_0_317<=Wgt_0_317; w_0_318<=Wgt_0_318; w_0_319<=Wgt_0_319; w_0_320<=Wgt_0_320; w_0_321<=Wgt_0_321; w_0_322<=Wgt_0_322; w_0_323<=Wgt_0_323; w_0_324<=Wgt_0_324; w_0_325<=Wgt_0_325; w_0_326<=Wgt_0_326; w_0_327<=Wgt_0_327; w_0_328<=Wgt_0_328; w_0_329<=Wgt_0_329; w_0_330<=Wgt_0_330; w_0_331<=Wgt_0_331; w_0_332<=Wgt_0_332; w_0_333<=Wgt_0_333; w_0_334<=Wgt_0_334; w_0_335<=Wgt_0_335; w_0_336<=Wgt_0_336; w_0_337<=Wgt_0_337; w_0_338<=Wgt_0_338; w_0_339<=Wgt_0_339; w_0_340<=Wgt_0_340; w_0_341<=Wgt_0_341; w_0_342<=Wgt_0_342; w_0_343<=Wgt_0_343; w_0_344<=Wgt_0_344; w_0_345<=Wgt_0_345; w_0_346<=Wgt_0_346; w_0_347<=Wgt_0_347; w_0_348<=Wgt_0_348; w_0_349<=Wgt_0_349; w_0_350<=Wgt_0_350; w_0_351<=Wgt_0_351; w_0_352<=Wgt_0_352; w_0_353<=Wgt_0_353; w_0_354<=Wgt_0_354; w_0_355<=Wgt_0_355; w_0_356<=Wgt_0_356; w_0_357<=Wgt_0_357; w_0_358<=Wgt_0_358; w_0_359<=Wgt_0_359; w_0_360<=Wgt_0_360; w_0_361<=Wgt_0_361; w_0_362<=Wgt_0_362; w_0_363<=Wgt_0_363; w_0_364<=Wgt_0_364; w_0_365<=Wgt_0_365; w_0_366<=Wgt_0_366; w_0_367<=Wgt_0_367; w_0_368<=Wgt_0_368; w_0_369<=Wgt_0_369; w_0_370<=Wgt_0_370; w_0_371<=Wgt_0_371; w_0_372<=Wgt_0_372; w_0_373<=Wgt_0_373; w_0_374<=Wgt_0_374; w_0_375<=Wgt_0_375; w_0_376<=Wgt_0_376; w_0_377<=Wgt_0_377; w_0_378<=Wgt_0_378; w_0_379<=Wgt_0_379; w_0_380<=Wgt_0_380; w_0_381<=Wgt_0_381; w_0_382<=Wgt_0_382; w_0_383<=Wgt_0_383; w_0_384<=Wgt_0_384; w_0_385<=Wgt_0_385; w_0_386<=Wgt_0_386; w_0_387<=Wgt_0_387; w_0_388<=Wgt_0_388; w_0_389<=Wgt_0_389; w_0_390<=Wgt_0_390; w_0_391<=Wgt_0_391; w_0_392<=Wgt_0_392; w_0_393<=Wgt_0_393; w_0_394<=Wgt_0_394; w_0_395<=Wgt_0_395; w_0_396<=Wgt_0_396; w_0_397<=Wgt_0_397; w_0_398<=Wgt_0_398; w_0_399<=Wgt_0_399; w_0_400<=Wgt_0_400; w_0_401<=Wgt_0_401; w_0_402<=Wgt_0_402; w_0_403<=Wgt_0_403; w_0_404<=Wgt_0_404; w_0_405<=Wgt_0_405; w_0_406<=Wgt_0_406; w_0_407<=Wgt_0_407; w_0_408<=Wgt_0_408; w_0_409<=Wgt_0_409; w_0_410<=Wgt_0_410; w_0_411<=Wgt_0_411; w_0_412<=Wgt_0_412; w_0_413<=Wgt_0_413; w_0_414<=Wgt_0_414; w_0_415<=Wgt_0_415; w_0_416<=Wgt_0_416; w_0_417<=Wgt_0_417; w_0_418<=Wgt_0_418; w_0_419<=Wgt_0_419; w_0_420<=Wgt_0_420; w_0_421<=Wgt_0_421; w_0_422<=Wgt_0_422; w_0_423<=Wgt_0_423; w_0_424<=Wgt_0_424; w_0_425<=Wgt_0_425; w_0_426<=Wgt_0_426; w_0_427<=Wgt_0_427; w_0_428<=Wgt_0_428; w_0_429<=Wgt_0_429; w_0_430<=Wgt_0_430; w_0_431<=Wgt_0_431; w_0_432<=Wgt_0_432; w_0_433<=Wgt_0_433; w_0_434<=Wgt_0_434; w_0_435<=Wgt_0_435; w_0_436<=Wgt_0_436; w_0_437<=Wgt_0_437; w_0_438<=Wgt_0_438; w_0_439<=Wgt_0_439; w_0_440<=Wgt_0_440; w_0_441<=Wgt_0_441; w_0_442<=Wgt_0_442; w_0_443<=Wgt_0_443; w_0_444<=Wgt_0_444; w_0_445<=Wgt_0_445; w_0_446<=Wgt_0_446; w_0_447<=Wgt_0_447; w_0_448<=Wgt_0_448; w_0_449<=Wgt_0_449; w_0_450<=Wgt_0_450; w_0_451<=Wgt_0_451; w_0_452<=Wgt_0_452; w_0_453<=Wgt_0_453; w_0_454<=Wgt_0_454; w_0_455<=Wgt_0_455; w_0_456<=Wgt_0_456; w_0_457<=Wgt_0_457; w_0_458<=Wgt_0_458; w_0_459<=Wgt_0_459; w_0_460<=Wgt_0_460; w_0_461<=Wgt_0_461; w_0_462<=Wgt_0_462; w_0_463<=Wgt_0_463; w_0_464<=Wgt_0_464; w_0_465<=Wgt_0_465; w_0_466<=Wgt_0_466; w_0_467<=Wgt_0_467; w_0_468<=Wgt_0_468; w_0_469<=Wgt_0_469; w_0_470<=Wgt_0_470; w_0_471<=Wgt_0_471; w_0_472<=Wgt_0_472; w_0_473<=Wgt_0_473; w_0_474<=Wgt_0_474; w_0_475<=Wgt_0_475; w_0_476<=Wgt_0_476; w_0_477<=Wgt_0_477; w_0_478<=Wgt_0_478; w_0_479<=Wgt_0_479; w_0_480<=Wgt_0_480; w_0_481<=Wgt_0_481; w_0_482<=Wgt_0_482; w_0_483<=Wgt_0_483; w_0_484<=Wgt_0_484; w_0_485<=Wgt_0_485; w_0_486<=Wgt_0_486; w_0_487<=Wgt_0_487; w_0_488<=Wgt_0_488; w_0_489<=Wgt_0_489; w_0_490<=Wgt_0_490; w_0_491<=Wgt_0_491; w_0_492<=Wgt_0_492; w_0_493<=Wgt_0_493; w_0_494<=Wgt_0_494; w_0_495<=Wgt_0_495; w_0_496<=Wgt_0_496; w_0_497<=Wgt_0_497; w_0_498<=Wgt_0_498; w_0_499<=Wgt_0_499; w_0_500<=Wgt_0_500; w_0_501<=Wgt_0_501; w_0_502<=Wgt_0_502; w_0_503<=Wgt_0_503; w_0_504<=Wgt_0_504; w_0_505<=Wgt_0_505; w_0_506<=Wgt_0_506; w_0_507<=Wgt_0_507; w_0_508<=Wgt_0_508; w_0_509<=Wgt_0_509; w_0_510<=Wgt_0_510; w_0_511<=Wgt_0_511; w_0_512<=Wgt_0_512; w_0_513<=Wgt_0_513; w_0_514<=Wgt_0_514; w_0_515<=Wgt_0_515; w_0_516<=Wgt_0_516; w_0_517<=Wgt_0_517; w_0_518<=Wgt_0_518; w_0_519<=Wgt_0_519; w_0_520<=Wgt_0_520; w_0_521<=Wgt_0_521; w_0_522<=Wgt_0_522; w_0_523<=Wgt_0_523; w_0_524<=Wgt_0_524; w_0_525<=Wgt_0_525; w_0_526<=Wgt_0_526; w_0_527<=Wgt_0_527; w_0_528<=Wgt_0_528; w_0_529<=Wgt_0_529; w_0_530<=Wgt_0_530; w_0_531<=Wgt_0_531; w_0_532<=Wgt_0_532; w_0_533<=Wgt_0_533; w_0_534<=Wgt_0_534; w_0_535<=Wgt_0_535; w_0_536<=Wgt_0_536; w_0_537<=Wgt_0_537; w_0_538<=Wgt_0_538; w_0_539<=Wgt_0_539; w_0_540<=Wgt_0_540; w_0_541<=Wgt_0_541; w_0_542<=Wgt_0_542; w_0_543<=Wgt_0_543; w_0_544<=Wgt_0_544; w_0_545<=Wgt_0_545; w_0_546<=Wgt_0_546; w_0_547<=Wgt_0_547; w_0_548<=Wgt_0_548; w_0_549<=Wgt_0_549; w_0_550<=Wgt_0_550; w_0_551<=Wgt_0_551; w_0_552<=Wgt_0_552; w_0_553<=Wgt_0_553; w_0_554<=Wgt_0_554; w_0_555<=Wgt_0_555; w_0_556<=Wgt_0_556; w_0_557<=Wgt_0_557; w_0_558<=Wgt_0_558; w_0_559<=Wgt_0_559; w_0_560<=Wgt_0_560; w_0_561<=Wgt_0_561; w_0_562<=Wgt_0_562; w_0_563<=Wgt_0_563; w_0_564<=Wgt_0_564; w_0_565<=Wgt_0_565; w_0_566<=Wgt_0_566; w_0_567<=Wgt_0_567; w_0_568<=Wgt_0_568; w_0_569<=Wgt_0_569; w_0_570<=Wgt_0_570; w_0_571<=Wgt_0_571; w_0_572<=Wgt_0_572; w_0_573<=Wgt_0_573; w_0_574<=Wgt_0_574; w_0_575<=Wgt_0_575; w_0_576<=Wgt_0_576; w_0_577<=Wgt_0_577; w_0_578<=Wgt_0_578; w_0_579<=Wgt_0_579; w_0_580<=Wgt_0_580; w_0_581<=Wgt_0_581; w_0_582<=Wgt_0_582; w_0_583<=Wgt_0_583; w_0_584<=Wgt_0_584; w_0_585<=Wgt_0_585; w_0_586<=Wgt_0_586; w_0_587<=Wgt_0_587; w_0_588<=Wgt_0_588; w_0_589<=Wgt_0_589; w_0_590<=Wgt_0_590; w_0_591<=Wgt_0_591; w_0_592<=Wgt_0_592; w_0_593<=Wgt_0_593; w_0_594<=Wgt_0_594; w_0_595<=Wgt_0_595; w_0_596<=Wgt_0_596; w_0_597<=Wgt_0_597; w_0_598<=Wgt_0_598; w_0_599<=Wgt_0_599; w_0_600<=Wgt_0_600; w_0_601<=Wgt_0_601; w_0_602<=Wgt_0_602; w_0_603<=Wgt_0_603; w_0_604<=Wgt_0_604; w_0_605<=Wgt_0_605; w_0_606<=Wgt_0_606; w_0_607<=Wgt_0_607; w_0_608<=Wgt_0_608; w_0_609<=Wgt_0_609; w_0_610<=Wgt_0_610; w_0_611<=Wgt_0_611; w_0_612<=Wgt_0_612; w_0_613<=Wgt_0_613; w_0_614<=Wgt_0_614; w_0_615<=Wgt_0_615; w_0_616<=Wgt_0_616; w_0_617<=Wgt_0_617; w_0_618<=Wgt_0_618; w_0_619<=Wgt_0_619; w_0_620<=Wgt_0_620; w_0_621<=Wgt_0_621; w_0_622<=Wgt_0_622; w_0_623<=Wgt_0_623; w_0_624<=Wgt_0_624; w_0_625<=Wgt_0_625; w_0_626<=Wgt_0_626; w_0_627<=Wgt_0_627; w_0_628<=Wgt_0_628; w_0_629<=Wgt_0_629; w_0_630<=Wgt_0_630; w_0_631<=Wgt_0_631; w_0_632<=Wgt_0_632; w_0_633<=Wgt_0_633; w_0_634<=Wgt_0_634; w_0_635<=Wgt_0_635; w_0_636<=Wgt_0_636; w_0_637<=Wgt_0_637; w_0_638<=Wgt_0_638; w_0_639<=Wgt_0_639; w_0_640<=Wgt_0_640; w_0_641<=Wgt_0_641; w_0_642<=Wgt_0_642; w_0_643<=Wgt_0_643; w_0_644<=Wgt_0_644; w_0_645<=Wgt_0_645; w_0_646<=Wgt_0_646; w_0_647<=Wgt_0_647; w_0_648<=Wgt_0_648; w_0_649<=Wgt_0_649; w_0_650<=Wgt_0_650; w_0_651<=Wgt_0_651; w_0_652<=Wgt_0_652; w_0_653<=Wgt_0_653; w_0_654<=Wgt_0_654; w_0_655<=Wgt_0_655; w_0_656<=Wgt_0_656; w_0_657<=Wgt_0_657; w_0_658<=Wgt_0_658; w_0_659<=Wgt_0_659; w_0_660<=Wgt_0_660; w_0_661<=Wgt_0_661; w_0_662<=Wgt_0_662; w_0_663<=Wgt_0_663; w_0_664<=Wgt_0_664; w_0_665<=Wgt_0_665; w_0_666<=Wgt_0_666; w_0_667<=Wgt_0_667; w_0_668<=Wgt_0_668; w_0_669<=Wgt_0_669; w_0_670<=Wgt_0_670; w_0_671<=Wgt_0_671; w_0_672<=Wgt_0_672; w_0_673<=Wgt_0_673; w_0_674<=Wgt_0_674; w_0_675<=Wgt_0_675; w_0_676<=Wgt_0_676; w_0_677<=Wgt_0_677; w_0_678<=Wgt_0_678; w_0_679<=Wgt_0_679; w_0_680<=Wgt_0_680; w_0_681<=Wgt_0_681; w_0_682<=Wgt_0_682; w_0_683<=Wgt_0_683; w_0_684<=Wgt_0_684; w_0_685<=Wgt_0_685; w_0_686<=Wgt_0_686; w_0_687<=Wgt_0_687; w_0_688<=Wgt_0_688; w_0_689<=Wgt_0_689; w_0_690<=Wgt_0_690; w_0_691<=Wgt_0_691; w_0_692<=Wgt_0_692; w_0_693<=Wgt_0_693; w_0_694<=Wgt_0_694; w_0_695<=Wgt_0_695; w_0_696<=Wgt_0_696; w_0_697<=Wgt_0_697; w_0_698<=Wgt_0_698; w_0_699<=Wgt_0_699; w_0_700<=Wgt_0_700; w_0_701<=Wgt_0_701; w_0_702<=Wgt_0_702; w_0_703<=Wgt_0_703; w_0_704<=Wgt_0_704; w_0_705<=Wgt_0_705; w_0_706<=Wgt_0_706; w_0_707<=Wgt_0_707; w_0_708<=Wgt_0_708; w_0_709<=Wgt_0_709; w_0_710<=Wgt_0_710; w_0_711<=Wgt_0_711; w_0_712<=Wgt_0_712; w_0_713<=Wgt_0_713; w_0_714<=Wgt_0_714; w_0_715<=Wgt_0_715; w_0_716<=Wgt_0_716; w_0_717<=Wgt_0_717; w_0_718<=Wgt_0_718; w_0_719<=Wgt_0_719; w_0_720<=Wgt_0_720; w_0_721<=Wgt_0_721; w_0_722<=Wgt_0_722; w_0_723<=Wgt_0_723; w_0_724<=Wgt_0_724; w_0_725<=Wgt_0_725; w_0_726<=Wgt_0_726; w_0_727<=Wgt_0_727; w_0_728<=Wgt_0_728; w_0_729<=Wgt_0_729; w_0_730<=Wgt_0_730; w_0_731<=Wgt_0_731; w_0_732<=Wgt_0_732; w_0_733<=Wgt_0_733; w_0_734<=Wgt_0_734; w_0_735<=Wgt_0_735; w_0_736<=Wgt_0_736; w_0_737<=Wgt_0_737; w_0_738<=Wgt_0_738; w_0_739<=Wgt_0_739; w_0_740<=Wgt_0_740; w_0_741<=Wgt_0_741; w_0_742<=Wgt_0_742; w_0_743<=Wgt_0_743; w_0_744<=Wgt_0_744; w_0_745<=Wgt_0_745; w_0_746<=Wgt_0_746; w_0_747<=Wgt_0_747; w_0_748<=Wgt_0_748; w_0_749<=Wgt_0_749; w_0_750<=Wgt_0_750; w_0_751<=Wgt_0_751; w_0_752<=Wgt_0_752; w_0_753<=Wgt_0_753; w_0_754<=Wgt_0_754; w_0_755<=Wgt_0_755; w_0_756<=Wgt_0_756; w_0_757<=Wgt_0_757; w_0_758<=Wgt_0_758; w_0_759<=Wgt_0_759; w_0_760<=Wgt_0_760; w_0_761<=Wgt_0_761; w_0_762<=Wgt_0_762; w_0_763<=Wgt_0_763; w_0_764<=Wgt_0_764; w_0_765<=Wgt_0_765; w_0_766<=Wgt_0_766; w_0_767<=Wgt_0_767; w_0_768<=Wgt_0_768; w_0_769<=Wgt_0_769; w_0_770<=Wgt_0_770; w_0_771<=Wgt_0_771; w_0_772<=Wgt_0_772; w_0_773<=Wgt_0_773; w_0_774<=Wgt_0_774; w_0_775<=Wgt_0_775; w_0_776<=Wgt_0_776; w_0_777<=Wgt_0_777; w_0_778<=Wgt_0_778; w_0_779<=Wgt_0_779; w_0_780<=Wgt_0_780; w_0_781<=Wgt_0_781; w_0_782<=Wgt_0_782; w_0_783<=Wgt_0_783; w_0_784<=Wgt_0_784; 
					w_1_0<=Wgt_1_0; w_1_1<=Wgt_1_1; w_1_2<=Wgt_1_2; w_1_3<=Wgt_1_3; w_1_4<=Wgt_1_4; w_1_5<=Wgt_1_5; w_1_6<=Wgt_1_6; w_1_7<=Wgt_1_7; w_1_8<=Wgt_1_8; w_1_9<=Wgt_1_9; w_1_10<=Wgt_1_10; w_1_11<=Wgt_1_11; w_1_12<=Wgt_1_12; w_1_13<=Wgt_1_13; w_1_14<=Wgt_1_14; w_1_15<=Wgt_1_15; w_1_16<=Wgt_1_16; w_1_17<=Wgt_1_17; w_1_18<=Wgt_1_18; w_1_19<=Wgt_1_19; w_1_20<=Wgt_1_20; w_1_21<=Wgt_1_21; w_1_22<=Wgt_1_22; w_1_23<=Wgt_1_23; w_1_24<=Wgt_1_24; w_1_25<=Wgt_1_25; w_1_26<=Wgt_1_26; w_1_27<=Wgt_1_27; w_1_28<=Wgt_1_28; w_1_29<=Wgt_1_29; w_1_30<=Wgt_1_30; w_1_31<=Wgt_1_31; w_1_32<=Wgt_1_32; w_1_33<=Wgt_1_33; w_1_34<=Wgt_1_34; w_1_35<=Wgt_1_35; w_1_36<=Wgt_1_36; w_1_37<=Wgt_1_37; w_1_38<=Wgt_1_38; w_1_39<=Wgt_1_39; w_1_40<=Wgt_1_40; w_1_41<=Wgt_1_41; w_1_42<=Wgt_1_42; w_1_43<=Wgt_1_43; w_1_44<=Wgt_1_44; w_1_45<=Wgt_1_45; w_1_46<=Wgt_1_46; w_1_47<=Wgt_1_47; w_1_48<=Wgt_1_48; w_1_49<=Wgt_1_49; w_1_50<=Wgt_1_50; w_1_51<=Wgt_1_51; w_1_52<=Wgt_1_52; w_1_53<=Wgt_1_53; w_1_54<=Wgt_1_54; w_1_55<=Wgt_1_55; w_1_56<=Wgt_1_56; w_1_57<=Wgt_1_57; w_1_58<=Wgt_1_58; w_1_59<=Wgt_1_59; w_1_60<=Wgt_1_60; w_1_61<=Wgt_1_61; w_1_62<=Wgt_1_62; w_1_63<=Wgt_1_63; w_1_64<=Wgt_1_64; w_1_65<=Wgt_1_65; w_1_66<=Wgt_1_66; w_1_67<=Wgt_1_67; w_1_68<=Wgt_1_68; w_1_69<=Wgt_1_69; w_1_70<=Wgt_1_70; w_1_71<=Wgt_1_71; w_1_72<=Wgt_1_72; w_1_73<=Wgt_1_73; w_1_74<=Wgt_1_74; w_1_75<=Wgt_1_75; w_1_76<=Wgt_1_76; w_1_77<=Wgt_1_77; w_1_78<=Wgt_1_78; w_1_79<=Wgt_1_79; w_1_80<=Wgt_1_80; w_1_81<=Wgt_1_81; w_1_82<=Wgt_1_82; w_1_83<=Wgt_1_83; w_1_84<=Wgt_1_84; w_1_85<=Wgt_1_85; w_1_86<=Wgt_1_86; w_1_87<=Wgt_1_87; w_1_88<=Wgt_1_88; w_1_89<=Wgt_1_89; w_1_90<=Wgt_1_90; w_1_91<=Wgt_1_91; w_1_92<=Wgt_1_92; w_1_93<=Wgt_1_93; w_1_94<=Wgt_1_94; w_1_95<=Wgt_1_95; w_1_96<=Wgt_1_96; w_1_97<=Wgt_1_97; w_1_98<=Wgt_1_98; w_1_99<=Wgt_1_99; w_1_100<=Wgt_1_100; w_1_101<=Wgt_1_101; w_1_102<=Wgt_1_102; w_1_103<=Wgt_1_103; w_1_104<=Wgt_1_104; w_1_105<=Wgt_1_105; w_1_106<=Wgt_1_106; w_1_107<=Wgt_1_107; w_1_108<=Wgt_1_108; w_1_109<=Wgt_1_109; w_1_110<=Wgt_1_110; w_1_111<=Wgt_1_111; w_1_112<=Wgt_1_112; w_1_113<=Wgt_1_113; w_1_114<=Wgt_1_114; w_1_115<=Wgt_1_115; w_1_116<=Wgt_1_116; w_1_117<=Wgt_1_117; w_1_118<=Wgt_1_118; w_1_119<=Wgt_1_119; w_1_120<=Wgt_1_120; w_1_121<=Wgt_1_121; w_1_122<=Wgt_1_122; w_1_123<=Wgt_1_123; w_1_124<=Wgt_1_124; w_1_125<=Wgt_1_125; w_1_126<=Wgt_1_126; w_1_127<=Wgt_1_127; w_1_128<=Wgt_1_128; w_1_129<=Wgt_1_129; w_1_130<=Wgt_1_130; w_1_131<=Wgt_1_131; w_1_132<=Wgt_1_132; w_1_133<=Wgt_1_133; w_1_134<=Wgt_1_134; w_1_135<=Wgt_1_135; w_1_136<=Wgt_1_136; w_1_137<=Wgt_1_137; w_1_138<=Wgt_1_138; w_1_139<=Wgt_1_139; w_1_140<=Wgt_1_140; w_1_141<=Wgt_1_141; w_1_142<=Wgt_1_142; w_1_143<=Wgt_1_143; w_1_144<=Wgt_1_144; w_1_145<=Wgt_1_145; w_1_146<=Wgt_1_146; w_1_147<=Wgt_1_147; w_1_148<=Wgt_1_148; w_1_149<=Wgt_1_149; w_1_150<=Wgt_1_150; w_1_151<=Wgt_1_151; w_1_152<=Wgt_1_152; w_1_153<=Wgt_1_153; w_1_154<=Wgt_1_154; w_1_155<=Wgt_1_155; w_1_156<=Wgt_1_156; w_1_157<=Wgt_1_157; w_1_158<=Wgt_1_158; w_1_159<=Wgt_1_159; w_1_160<=Wgt_1_160; w_1_161<=Wgt_1_161; w_1_162<=Wgt_1_162; w_1_163<=Wgt_1_163; w_1_164<=Wgt_1_164; w_1_165<=Wgt_1_165; w_1_166<=Wgt_1_166; w_1_167<=Wgt_1_167; w_1_168<=Wgt_1_168; w_1_169<=Wgt_1_169; w_1_170<=Wgt_1_170; w_1_171<=Wgt_1_171; w_1_172<=Wgt_1_172; w_1_173<=Wgt_1_173; w_1_174<=Wgt_1_174; w_1_175<=Wgt_1_175; w_1_176<=Wgt_1_176; w_1_177<=Wgt_1_177; w_1_178<=Wgt_1_178; w_1_179<=Wgt_1_179; w_1_180<=Wgt_1_180; w_1_181<=Wgt_1_181; w_1_182<=Wgt_1_182; w_1_183<=Wgt_1_183; w_1_184<=Wgt_1_184; w_1_185<=Wgt_1_185; w_1_186<=Wgt_1_186; w_1_187<=Wgt_1_187; w_1_188<=Wgt_1_188; w_1_189<=Wgt_1_189; w_1_190<=Wgt_1_190; w_1_191<=Wgt_1_191; w_1_192<=Wgt_1_192; w_1_193<=Wgt_1_193; w_1_194<=Wgt_1_194; w_1_195<=Wgt_1_195; w_1_196<=Wgt_1_196; w_1_197<=Wgt_1_197; w_1_198<=Wgt_1_198; w_1_199<=Wgt_1_199; w_1_200<=Wgt_1_200; w_1_201<=Wgt_1_201; w_1_202<=Wgt_1_202; w_1_203<=Wgt_1_203; w_1_204<=Wgt_1_204; w_1_205<=Wgt_1_205; w_1_206<=Wgt_1_206; w_1_207<=Wgt_1_207; w_1_208<=Wgt_1_208; w_1_209<=Wgt_1_209; w_1_210<=Wgt_1_210; w_1_211<=Wgt_1_211; w_1_212<=Wgt_1_212; w_1_213<=Wgt_1_213; w_1_214<=Wgt_1_214; w_1_215<=Wgt_1_215; w_1_216<=Wgt_1_216; w_1_217<=Wgt_1_217; w_1_218<=Wgt_1_218; w_1_219<=Wgt_1_219; w_1_220<=Wgt_1_220; w_1_221<=Wgt_1_221; w_1_222<=Wgt_1_222; w_1_223<=Wgt_1_223; w_1_224<=Wgt_1_224; w_1_225<=Wgt_1_225; w_1_226<=Wgt_1_226; w_1_227<=Wgt_1_227; w_1_228<=Wgt_1_228; w_1_229<=Wgt_1_229; w_1_230<=Wgt_1_230; w_1_231<=Wgt_1_231; w_1_232<=Wgt_1_232; w_1_233<=Wgt_1_233; w_1_234<=Wgt_1_234; w_1_235<=Wgt_1_235; w_1_236<=Wgt_1_236; w_1_237<=Wgt_1_237; w_1_238<=Wgt_1_238; w_1_239<=Wgt_1_239; w_1_240<=Wgt_1_240; w_1_241<=Wgt_1_241; w_1_242<=Wgt_1_242; w_1_243<=Wgt_1_243; w_1_244<=Wgt_1_244; w_1_245<=Wgt_1_245; w_1_246<=Wgt_1_246; w_1_247<=Wgt_1_247; w_1_248<=Wgt_1_248; w_1_249<=Wgt_1_249; w_1_250<=Wgt_1_250; w_1_251<=Wgt_1_251; w_1_252<=Wgt_1_252; w_1_253<=Wgt_1_253; w_1_254<=Wgt_1_254; w_1_255<=Wgt_1_255; w_1_256<=Wgt_1_256; w_1_257<=Wgt_1_257; w_1_258<=Wgt_1_258; w_1_259<=Wgt_1_259; w_1_260<=Wgt_1_260; w_1_261<=Wgt_1_261; w_1_262<=Wgt_1_262; w_1_263<=Wgt_1_263; w_1_264<=Wgt_1_264; w_1_265<=Wgt_1_265; w_1_266<=Wgt_1_266; w_1_267<=Wgt_1_267; w_1_268<=Wgt_1_268; w_1_269<=Wgt_1_269; w_1_270<=Wgt_1_270; w_1_271<=Wgt_1_271; w_1_272<=Wgt_1_272; w_1_273<=Wgt_1_273; w_1_274<=Wgt_1_274; w_1_275<=Wgt_1_275; w_1_276<=Wgt_1_276; w_1_277<=Wgt_1_277; w_1_278<=Wgt_1_278; w_1_279<=Wgt_1_279; w_1_280<=Wgt_1_280; w_1_281<=Wgt_1_281; w_1_282<=Wgt_1_282; w_1_283<=Wgt_1_283; w_1_284<=Wgt_1_284; w_1_285<=Wgt_1_285; w_1_286<=Wgt_1_286; w_1_287<=Wgt_1_287; w_1_288<=Wgt_1_288; w_1_289<=Wgt_1_289; w_1_290<=Wgt_1_290; w_1_291<=Wgt_1_291; w_1_292<=Wgt_1_292; w_1_293<=Wgt_1_293; w_1_294<=Wgt_1_294; w_1_295<=Wgt_1_295; w_1_296<=Wgt_1_296; w_1_297<=Wgt_1_297; w_1_298<=Wgt_1_298; w_1_299<=Wgt_1_299; w_1_300<=Wgt_1_300; w_1_301<=Wgt_1_301; w_1_302<=Wgt_1_302; w_1_303<=Wgt_1_303; w_1_304<=Wgt_1_304; w_1_305<=Wgt_1_305; w_1_306<=Wgt_1_306; w_1_307<=Wgt_1_307; w_1_308<=Wgt_1_308; w_1_309<=Wgt_1_309; w_1_310<=Wgt_1_310; w_1_311<=Wgt_1_311; w_1_312<=Wgt_1_312; w_1_313<=Wgt_1_313; w_1_314<=Wgt_1_314; w_1_315<=Wgt_1_315; w_1_316<=Wgt_1_316; w_1_317<=Wgt_1_317; w_1_318<=Wgt_1_318; w_1_319<=Wgt_1_319; w_1_320<=Wgt_1_320; w_1_321<=Wgt_1_321; w_1_322<=Wgt_1_322; w_1_323<=Wgt_1_323; w_1_324<=Wgt_1_324; w_1_325<=Wgt_1_325; w_1_326<=Wgt_1_326; w_1_327<=Wgt_1_327; w_1_328<=Wgt_1_328; w_1_329<=Wgt_1_329; w_1_330<=Wgt_1_330; w_1_331<=Wgt_1_331; w_1_332<=Wgt_1_332; w_1_333<=Wgt_1_333; w_1_334<=Wgt_1_334; w_1_335<=Wgt_1_335; w_1_336<=Wgt_1_336; w_1_337<=Wgt_1_337; w_1_338<=Wgt_1_338; w_1_339<=Wgt_1_339; w_1_340<=Wgt_1_340; w_1_341<=Wgt_1_341; w_1_342<=Wgt_1_342; w_1_343<=Wgt_1_343; w_1_344<=Wgt_1_344; w_1_345<=Wgt_1_345; w_1_346<=Wgt_1_346; w_1_347<=Wgt_1_347; w_1_348<=Wgt_1_348; w_1_349<=Wgt_1_349; w_1_350<=Wgt_1_350; w_1_351<=Wgt_1_351; w_1_352<=Wgt_1_352; w_1_353<=Wgt_1_353; w_1_354<=Wgt_1_354; w_1_355<=Wgt_1_355; w_1_356<=Wgt_1_356; w_1_357<=Wgt_1_357; w_1_358<=Wgt_1_358; w_1_359<=Wgt_1_359; w_1_360<=Wgt_1_360; w_1_361<=Wgt_1_361; w_1_362<=Wgt_1_362; w_1_363<=Wgt_1_363; w_1_364<=Wgt_1_364; w_1_365<=Wgt_1_365; w_1_366<=Wgt_1_366; w_1_367<=Wgt_1_367; w_1_368<=Wgt_1_368; w_1_369<=Wgt_1_369; w_1_370<=Wgt_1_370; w_1_371<=Wgt_1_371; w_1_372<=Wgt_1_372; w_1_373<=Wgt_1_373; w_1_374<=Wgt_1_374; w_1_375<=Wgt_1_375; w_1_376<=Wgt_1_376; w_1_377<=Wgt_1_377; w_1_378<=Wgt_1_378; w_1_379<=Wgt_1_379; w_1_380<=Wgt_1_380; w_1_381<=Wgt_1_381; w_1_382<=Wgt_1_382; w_1_383<=Wgt_1_383; w_1_384<=Wgt_1_384; w_1_385<=Wgt_1_385; w_1_386<=Wgt_1_386; w_1_387<=Wgt_1_387; w_1_388<=Wgt_1_388; w_1_389<=Wgt_1_389; w_1_390<=Wgt_1_390; w_1_391<=Wgt_1_391; w_1_392<=Wgt_1_392; w_1_393<=Wgt_1_393; w_1_394<=Wgt_1_394; w_1_395<=Wgt_1_395; w_1_396<=Wgt_1_396; w_1_397<=Wgt_1_397; w_1_398<=Wgt_1_398; w_1_399<=Wgt_1_399; w_1_400<=Wgt_1_400; w_1_401<=Wgt_1_401; w_1_402<=Wgt_1_402; w_1_403<=Wgt_1_403; w_1_404<=Wgt_1_404; w_1_405<=Wgt_1_405; w_1_406<=Wgt_1_406; w_1_407<=Wgt_1_407; w_1_408<=Wgt_1_408; w_1_409<=Wgt_1_409; w_1_410<=Wgt_1_410; w_1_411<=Wgt_1_411; w_1_412<=Wgt_1_412; w_1_413<=Wgt_1_413; w_1_414<=Wgt_1_414; w_1_415<=Wgt_1_415; w_1_416<=Wgt_1_416; w_1_417<=Wgt_1_417; w_1_418<=Wgt_1_418; w_1_419<=Wgt_1_419; w_1_420<=Wgt_1_420; w_1_421<=Wgt_1_421; w_1_422<=Wgt_1_422; w_1_423<=Wgt_1_423; w_1_424<=Wgt_1_424; w_1_425<=Wgt_1_425; w_1_426<=Wgt_1_426; w_1_427<=Wgt_1_427; w_1_428<=Wgt_1_428; w_1_429<=Wgt_1_429; w_1_430<=Wgt_1_430; w_1_431<=Wgt_1_431; w_1_432<=Wgt_1_432; w_1_433<=Wgt_1_433; w_1_434<=Wgt_1_434; w_1_435<=Wgt_1_435; w_1_436<=Wgt_1_436; w_1_437<=Wgt_1_437; w_1_438<=Wgt_1_438; w_1_439<=Wgt_1_439; w_1_440<=Wgt_1_440; w_1_441<=Wgt_1_441; w_1_442<=Wgt_1_442; w_1_443<=Wgt_1_443; w_1_444<=Wgt_1_444; w_1_445<=Wgt_1_445; w_1_446<=Wgt_1_446; w_1_447<=Wgt_1_447; w_1_448<=Wgt_1_448; w_1_449<=Wgt_1_449; w_1_450<=Wgt_1_450; w_1_451<=Wgt_1_451; w_1_452<=Wgt_1_452; w_1_453<=Wgt_1_453; w_1_454<=Wgt_1_454; w_1_455<=Wgt_1_455; w_1_456<=Wgt_1_456; w_1_457<=Wgt_1_457; w_1_458<=Wgt_1_458; w_1_459<=Wgt_1_459; w_1_460<=Wgt_1_460; w_1_461<=Wgt_1_461; w_1_462<=Wgt_1_462; w_1_463<=Wgt_1_463; w_1_464<=Wgt_1_464; w_1_465<=Wgt_1_465; w_1_466<=Wgt_1_466; w_1_467<=Wgt_1_467; w_1_468<=Wgt_1_468; w_1_469<=Wgt_1_469; w_1_470<=Wgt_1_470; w_1_471<=Wgt_1_471; w_1_472<=Wgt_1_472; w_1_473<=Wgt_1_473; w_1_474<=Wgt_1_474; w_1_475<=Wgt_1_475; w_1_476<=Wgt_1_476; w_1_477<=Wgt_1_477; w_1_478<=Wgt_1_478; w_1_479<=Wgt_1_479; w_1_480<=Wgt_1_480; w_1_481<=Wgt_1_481; w_1_482<=Wgt_1_482; w_1_483<=Wgt_1_483; w_1_484<=Wgt_1_484; w_1_485<=Wgt_1_485; w_1_486<=Wgt_1_486; w_1_487<=Wgt_1_487; w_1_488<=Wgt_1_488; w_1_489<=Wgt_1_489; w_1_490<=Wgt_1_490; w_1_491<=Wgt_1_491; w_1_492<=Wgt_1_492; w_1_493<=Wgt_1_493; w_1_494<=Wgt_1_494; w_1_495<=Wgt_1_495; w_1_496<=Wgt_1_496; w_1_497<=Wgt_1_497; w_1_498<=Wgt_1_498; w_1_499<=Wgt_1_499; w_1_500<=Wgt_1_500; w_1_501<=Wgt_1_501; w_1_502<=Wgt_1_502; w_1_503<=Wgt_1_503; w_1_504<=Wgt_1_504; w_1_505<=Wgt_1_505; w_1_506<=Wgt_1_506; w_1_507<=Wgt_1_507; w_1_508<=Wgt_1_508; w_1_509<=Wgt_1_509; w_1_510<=Wgt_1_510; w_1_511<=Wgt_1_511; w_1_512<=Wgt_1_512; w_1_513<=Wgt_1_513; w_1_514<=Wgt_1_514; w_1_515<=Wgt_1_515; w_1_516<=Wgt_1_516; w_1_517<=Wgt_1_517; w_1_518<=Wgt_1_518; w_1_519<=Wgt_1_519; w_1_520<=Wgt_1_520; w_1_521<=Wgt_1_521; w_1_522<=Wgt_1_522; w_1_523<=Wgt_1_523; w_1_524<=Wgt_1_524; w_1_525<=Wgt_1_525; w_1_526<=Wgt_1_526; w_1_527<=Wgt_1_527; w_1_528<=Wgt_1_528; w_1_529<=Wgt_1_529; w_1_530<=Wgt_1_530; w_1_531<=Wgt_1_531; w_1_532<=Wgt_1_532; w_1_533<=Wgt_1_533; w_1_534<=Wgt_1_534; w_1_535<=Wgt_1_535; w_1_536<=Wgt_1_536; w_1_537<=Wgt_1_537; w_1_538<=Wgt_1_538; w_1_539<=Wgt_1_539; w_1_540<=Wgt_1_540; w_1_541<=Wgt_1_541; w_1_542<=Wgt_1_542; w_1_543<=Wgt_1_543; w_1_544<=Wgt_1_544; w_1_545<=Wgt_1_545; w_1_546<=Wgt_1_546; w_1_547<=Wgt_1_547; w_1_548<=Wgt_1_548; w_1_549<=Wgt_1_549; w_1_550<=Wgt_1_550; w_1_551<=Wgt_1_551; w_1_552<=Wgt_1_552; w_1_553<=Wgt_1_553; w_1_554<=Wgt_1_554; w_1_555<=Wgt_1_555; w_1_556<=Wgt_1_556; w_1_557<=Wgt_1_557; w_1_558<=Wgt_1_558; w_1_559<=Wgt_1_559; w_1_560<=Wgt_1_560; w_1_561<=Wgt_1_561; w_1_562<=Wgt_1_562; w_1_563<=Wgt_1_563; w_1_564<=Wgt_1_564; w_1_565<=Wgt_1_565; w_1_566<=Wgt_1_566; w_1_567<=Wgt_1_567; w_1_568<=Wgt_1_568; w_1_569<=Wgt_1_569; w_1_570<=Wgt_1_570; w_1_571<=Wgt_1_571; w_1_572<=Wgt_1_572; w_1_573<=Wgt_1_573; w_1_574<=Wgt_1_574; w_1_575<=Wgt_1_575; w_1_576<=Wgt_1_576; w_1_577<=Wgt_1_577; w_1_578<=Wgt_1_578; w_1_579<=Wgt_1_579; w_1_580<=Wgt_1_580; w_1_581<=Wgt_1_581; w_1_582<=Wgt_1_582; w_1_583<=Wgt_1_583; w_1_584<=Wgt_1_584; w_1_585<=Wgt_1_585; w_1_586<=Wgt_1_586; w_1_587<=Wgt_1_587; w_1_588<=Wgt_1_588; w_1_589<=Wgt_1_589; w_1_590<=Wgt_1_590; w_1_591<=Wgt_1_591; w_1_592<=Wgt_1_592; w_1_593<=Wgt_1_593; w_1_594<=Wgt_1_594; w_1_595<=Wgt_1_595; w_1_596<=Wgt_1_596; w_1_597<=Wgt_1_597; w_1_598<=Wgt_1_598; w_1_599<=Wgt_1_599; w_1_600<=Wgt_1_600; w_1_601<=Wgt_1_601; w_1_602<=Wgt_1_602; w_1_603<=Wgt_1_603; w_1_604<=Wgt_1_604; w_1_605<=Wgt_1_605; w_1_606<=Wgt_1_606; w_1_607<=Wgt_1_607; w_1_608<=Wgt_1_608; w_1_609<=Wgt_1_609; w_1_610<=Wgt_1_610; w_1_611<=Wgt_1_611; w_1_612<=Wgt_1_612; w_1_613<=Wgt_1_613; w_1_614<=Wgt_1_614; w_1_615<=Wgt_1_615; w_1_616<=Wgt_1_616; w_1_617<=Wgt_1_617; w_1_618<=Wgt_1_618; w_1_619<=Wgt_1_619; w_1_620<=Wgt_1_620; w_1_621<=Wgt_1_621; w_1_622<=Wgt_1_622; w_1_623<=Wgt_1_623; w_1_624<=Wgt_1_624; w_1_625<=Wgt_1_625; w_1_626<=Wgt_1_626; w_1_627<=Wgt_1_627; w_1_628<=Wgt_1_628; w_1_629<=Wgt_1_629; w_1_630<=Wgt_1_630; w_1_631<=Wgt_1_631; w_1_632<=Wgt_1_632; w_1_633<=Wgt_1_633; w_1_634<=Wgt_1_634; w_1_635<=Wgt_1_635; w_1_636<=Wgt_1_636; w_1_637<=Wgt_1_637; w_1_638<=Wgt_1_638; w_1_639<=Wgt_1_639; w_1_640<=Wgt_1_640; w_1_641<=Wgt_1_641; w_1_642<=Wgt_1_642; w_1_643<=Wgt_1_643; w_1_644<=Wgt_1_644; w_1_645<=Wgt_1_645; w_1_646<=Wgt_1_646; w_1_647<=Wgt_1_647; w_1_648<=Wgt_1_648; w_1_649<=Wgt_1_649; w_1_650<=Wgt_1_650; w_1_651<=Wgt_1_651; w_1_652<=Wgt_1_652; w_1_653<=Wgt_1_653; w_1_654<=Wgt_1_654; w_1_655<=Wgt_1_655; w_1_656<=Wgt_1_656; w_1_657<=Wgt_1_657; w_1_658<=Wgt_1_658; w_1_659<=Wgt_1_659; w_1_660<=Wgt_1_660; w_1_661<=Wgt_1_661; w_1_662<=Wgt_1_662; w_1_663<=Wgt_1_663; w_1_664<=Wgt_1_664; w_1_665<=Wgt_1_665; w_1_666<=Wgt_1_666; w_1_667<=Wgt_1_667; w_1_668<=Wgt_1_668; w_1_669<=Wgt_1_669; w_1_670<=Wgt_1_670; w_1_671<=Wgt_1_671; w_1_672<=Wgt_1_672; w_1_673<=Wgt_1_673; w_1_674<=Wgt_1_674; w_1_675<=Wgt_1_675; w_1_676<=Wgt_1_676; w_1_677<=Wgt_1_677; w_1_678<=Wgt_1_678; w_1_679<=Wgt_1_679; w_1_680<=Wgt_1_680; w_1_681<=Wgt_1_681; w_1_682<=Wgt_1_682; w_1_683<=Wgt_1_683; w_1_684<=Wgt_1_684; w_1_685<=Wgt_1_685; w_1_686<=Wgt_1_686; w_1_687<=Wgt_1_687; w_1_688<=Wgt_1_688; w_1_689<=Wgt_1_689; w_1_690<=Wgt_1_690; w_1_691<=Wgt_1_691; w_1_692<=Wgt_1_692; w_1_693<=Wgt_1_693; w_1_694<=Wgt_1_694; w_1_695<=Wgt_1_695; w_1_696<=Wgt_1_696; w_1_697<=Wgt_1_697; w_1_698<=Wgt_1_698; w_1_699<=Wgt_1_699; w_1_700<=Wgt_1_700; w_1_701<=Wgt_1_701; w_1_702<=Wgt_1_702; w_1_703<=Wgt_1_703; w_1_704<=Wgt_1_704; w_1_705<=Wgt_1_705; w_1_706<=Wgt_1_706; w_1_707<=Wgt_1_707; w_1_708<=Wgt_1_708; w_1_709<=Wgt_1_709; w_1_710<=Wgt_1_710; w_1_711<=Wgt_1_711; w_1_712<=Wgt_1_712; w_1_713<=Wgt_1_713; w_1_714<=Wgt_1_714; w_1_715<=Wgt_1_715; w_1_716<=Wgt_1_716; w_1_717<=Wgt_1_717; w_1_718<=Wgt_1_718; w_1_719<=Wgt_1_719; w_1_720<=Wgt_1_720; w_1_721<=Wgt_1_721; w_1_722<=Wgt_1_722; w_1_723<=Wgt_1_723; w_1_724<=Wgt_1_724; w_1_725<=Wgt_1_725; w_1_726<=Wgt_1_726; w_1_727<=Wgt_1_727; w_1_728<=Wgt_1_728; w_1_729<=Wgt_1_729; w_1_730<=Wgt_1_730; w_1_731<=Wgt_1_731; w_1_732<=Wgt_1_732; w_1_733<=Wgt_1_733; w_1_734<=Wgt_1_734; w_1_735<=Wgt_1_735; w_1_736<=Wgt_1_736; w_1_737<=Wgt_1_737; w_1_738<=Wgt_1_738; w_1_739<=Wgt_1_739; w_1_740<=Wgt_1_740; w_1_741<=Wgt_1_741; w_1_742<=Wgt_1_742; w_1_743<=Wgt_1_743; w_1_744<=Wgt_1_744; w_1_745<=Wgt_1_745; w_1_746<=Wgt_1_746; w_1_747<=Wgt_1_747; w_1_748<=Wgt_1_748; w_1_749<=Wgt_1_749; w_1_750<=Wgt_1_750; w_1_751<=Wgt_1_751; w_1_752<=Wgt_1_752; w_1_753<=Wgt_1_753; w_1_754<=Wgt_1_754; w_1_755<=Wgt_1_755; w_1_756<=Wgt_1_756; w_1_757<=Wgt_1_757; w_1_758<=Wgt_1_758; w_1_759<=Wgt_1_759; w_1_760<=Wgt_1_760; w_1_761<=Wgt_1_761; w_1_762<=Wgt_1_762; w_1_763<=Wgt_1_763; w_1_764<=Wgt_1_764; w_1_765<=Wgt_1_765; w_1_766<=Wgt_1_766; w_1_767<=Wgt_1_767; w_1_768<=Wgt_1_768; w_1_769<=Wgt_1_769; w_1_770<=Wgt_1_770; w_1_771<=Wgt_1_771; w_1_772<=Wgt_1_772; w_1_773<=Wgt_1_773; w_1_774<=Wgt_1_774; w_1_775<=Wgt_1_775; w_1_776<=Wgt_1_776; w_1_777<=Wgt_1_777; w_1_778<=Wgt_1_778; w_1_779<=Wgt_1_779; w_1_780<=Wgt_1_780; w_1_781<=Wgt_1_781; w_1_782<=Wgt_1_782; w_1_783<=Wgt_1_783; w_1_784<=Wgt_1_784; 
					w_2_0<=Wgt_2_0; w_2_1<=Wgt_2_1; w_2_2<=Wgt_2_2; w_2_3<=Wgt_2_3; w_2_4<=Wgt_2_4; w_2_5<=Wgt_2_5; w_2_6<=Wgt_2_6; w_2_7<=Wgt_2_7; w_2_8<=Wgt_2_8; w_2_9<=Wgt_2_9; w_2_10<=Wgt_2_10; w_2_11<=Wgt_2_11; w_2_12<=Wgt_2_12; w_2_13<=Wgt_2_13; w_2_14<=Wgt_2_14; w_2_15<=Wgt_2_15; w_2_16<=Wgt_2_16; w_2_17<=Wgt_2_17; w_2_18<=Wgt_2_18; w_2_19<=Wgt_2_19; w_2_20<=Wgt_2_20; w_2_21<=Wgt_2_21; w_2_22<=Wgt_2_22; w_2_23<=Wgt_2_23; w_2_24<=Wgt_2_24; w_2_25<=Wgt_2_25; w_2_26<=Wgt_2_26; w_2_27<=Wgt_2_27; w_2_28<=Wgt_2_28; w_2_29<=Wgt_2_29; w_2_30<=Wgt_2_30; w_2_31<=Wgt_2_31; w_2_32<=Wgt_2_32; w_2_33<=Wgt_2_33; w_2_34<=Wgt_2_34; w_2_35<=Wgt_2_35; w_2_36<=Wgt_2_36; w_2_37<=Wgt_2_37; w_2_38<=Wgt_2_38; w_2_39<=Wgt_2_39; w_2_40<=Wgt_2_40; w_2_41<=Wgt_2_41; w_2_42<=Wgt_2_42; w_2_43<=Wgt_2_43; w_2_44<=Wgt_2_44; w_2_45<=Wgt_2_45; w_2_46<=Wgt_2_46; w_2_47<=Wgt_2_47; w_2_48<=Wgt_2_48; w_2_49<=Wgt_2_49; w_2_50<=Wgt_2_50; w_2_51<=Wgt_2_51; w_2_52<=Wgt_2_52; w_2_53<=Wgt_2_53; w_2_54<=Wgt_2_54; w_2_55<=Wgt_2_55; w_2_56<=Wgt_2_56; w_2_57<=Wgt_2_57; w_2_58<=Wgt_2_58; w_2_59<=Wgt_2_59; w_2_60<=Wgt_2_60; w_2_61<=Wgt_2_61; w_2_62<=Wgt_2_62; w_2_63<=Wgt_2_63; w_2_64<=Wgt_2_64; w_2_65<=Wgt_2_65; w_2_66<=Wgt_2_66; w_2_67<=Wgt_2_67; w_2_68<=Wgt_2_68; w_2_69<=Wgt_2_69; w_2_70<=Wgt_2_70; w_2_71<=Wgt_2_71; w_2_72<=Wgt_2_72; w_2_73<=Wgt_2_73; w_2_74<=Wgt_2_74; w_2_75<=Wgt_2_75; w_2_76<=Wgt_2_76; w_2_77<=Wgt_2_77; w_2_78<=Wgt_2_78; w_2_79<=Wgt_2_79; w_2_80<=Wgt_2_80; w_2_81<=Wgt_2_81; w_2_82<=Wgt_2_82; w_2_83<=Wgt_2_83; w_2_84<=Wgt_2_84; w_2_85<=Wgt_2_85; w_2_86<=Wgt_2_86; w_2_87<=Wgt_2_87; w_2_88<=Wgt_2_88; w_2_89<=Wgt_2_89; w_2_90<=Wgt_2_90; w_2_91<=Wgt_2_91; w_2_92<=Wgt_2_92; w_2_93<=Wgt_2_93; w_2_94<=Wgt_2_94; w_2_95<=Wgt_2_95; w_2_96<=Wgt_2_96; w_2_97<=Wgt_2_97; w_2_98<=Wgt_2_98; w_2_99<=Wgt_2_99; w_2_100<=Wgt_2_100; w_2_101<=Wgt_2_101; w_2_102<=Wgt_2_102; w_2_103<=Wgt_2_103; w_2_104<=Wgt_2_104; w_2_105<=Wgt_2_105; w_2_106<=Wgt_2_106; w_2_107<=Wgt_2_107; w_2_108<=Wgt_2_108; w_2_109<=Wgt_2_109; w_2_110<=Wgt_2_110; w_2_111<=Wgt_2_111; w_2_112<=Wgt_2_112; w_2_113<=Wgt_2_113; w_2_114<=Wgt_2_114; w_2_115<=Wgt_2_115; w_2_116<=Wgt_2_116; w_2_117<=Wgt_2_117; w_2_118<=Wgt_2_118; w_2_119<=Wgt_2_119; w_2_120<=Wgt_2_120; w_2_121<=Wgt_2_121; w_2_122<=Wgt_2_122; w_2_123<=Wgt_2_123; w_2_124<=Wgt_2_124; w_2_125<=Wgt_2_125; w_2_126<=Wgt_2_126; w_2_127<=Wgt_2_127; w_2_128<=Wgt_2_128; w_2_129<=Wgt_2_129; w_2_130<=Wgt_2_130; w_2_131<=Wgt_2_131; w_2_132<=Wgt_2_132; w_2_133<=Wgt_2_133; w_2_134<=Wgt_2_134; w_2_135<=Wgt_2_135; w_2_136<=Wgt_2_136; w_2_137<=Wgt_2_137; w_2_138<=Wgt_2_138; w_2_139<=Wgt_2_139; w_2_140<=Wgt_2_140; w_2_141<=Wgt_2_141; w_2_142<=Wgt_2_142; w_2_143<=Wgt_2_143; w_2_144<=Wgt_2_144; w_2_145<=Wgt_2_145; w_2_146<=Wgt_2_146; w_2_147<=Wgt_2_147; w_2_148<=Wgt_2_148; w_2_149<=Wgt_2_149; w_2_150<=Wgt_2_150; w_2_151<=Wgt_2_151; w_2_152<=Wgt_2_152; w_2_153<=Wgt_2_153; w_2_154<=Wgt_2_154; w_2_155<=Wgt_2_155; w_2_156<=Wgt_2_156; w_2_157<=Wgt_2_157; w_2_158<=Wgt_2_158; w_2_159<=Wgt_2_159; w_2_160<=Wgt_2_160; w_2_161<=Wgt_2_161; w_2_162<=Wgt_2_162; w_2_163<=Wgt_2_163; w_2_164<=Wgt_2_164; w_2_165<=Wgt_2_165; w_2_166<=Wgt_2_166; w_2_167<=Wgt_2_167; w_2_168<=Wgt_2_168; w_2_169<=Wgt_2_169; w_2_170<=Wgt_2_170; w_2_171<=Wgt_2_171; w_2_172<=Wgt_2_172; w_2_173<=Wgt_2_173; w_2_174<=Wgt_2_174; w_2_175<=Wgt_2_175; w_2_176<=Wgt_2_176; w_2_177<=Wgt_2_177; w_2_178<=Wgt_2_178; w_2_179<=Wgt_2_179; w_2_180<=Wgt_2_180; w_2_181<=Wgt_2_181; w_2_182<=Wgt_2_182; w_2_183<=Wgt_2_183; w_2_184<=Wgt_2_184; w_2_185<=Wgt_2_185; w_2_186<=Wgt_2_186; w_2_187<=Wgt_2_187; w_2_188<=Wgt_2_188; w_2_189<=Wgt_2_189; w_2_190<=Wgt_2_190; w_2_191<=Wgt_2_191; w_2_192<=Wgt_2_192; w_2_193<=Wgt_2_193; w_2_194<=Wgt_2_194; w_2_195<=Wgt_2_195; w_2_196<=Wgt_2_196; w_2_197<=Wgt_2_197; w_2_198<=Wgt_2_198; w_2_199<=Wgt_2_199; w_2_200<=Wgt_2_200; w_2_201<=Wgt_2_201; w_2_202<=Wgt_2_202; w_2_203<=Wgt_2_203; w_2_204<=Wgt_2_204; w_2_205<=Wgt_2_205; w_2_206<=Wgt_2_206; w_2_207<=Wgt_2_207; w_2_208<=Wgt_2_208; w_2_209<=Wgt_2_209; w_2_210<=Wgt_2_210; w_2_211<=Wgt_2_211; w_2_212<=Wgt_2_212; w_2_213<=Wgt_2_213; w_2_214<=Wgt_2_214; w_2_215<=Wgt_2_215; w_2_216<=Wgt_2_216; w_2_217<=Wgt_2_217; w_2_218<=Wgt_2_218; w_2_219<=Wgt_2_219; w_2_220<=Wgt_2_220; w_2_221<=Wgt_2_221; w_2_222<=Wgt_2_222; w_2_223<=Wgt_2_223; w_2_224<=Wgt_2_224; w_2_225<=Wgt_2_225; w_2_226<=Wgt_2_226; w_2_227<=Wgt_2_227; w_2_228<=Wgt_2_228; w_2_229<=Wgt_2_229; w_2_230<=Wgt_2_230; w_2_231<=Wgt_2_231; w_2_232<=Wgt_2_232; w_2_233<=Wgt_2_233; w_2_234<=Wgt_2_234; w_2_235<=Wgt_2_235; w_2_236<=Wgt_2_236; w_2_237<=Wgt_2_237; w_2_238<=Wgt_2_238; w_2_239<=Wgt_2_239; w_2_240<=Wgt_2_240; w_2_241<=Wgt_2_241; w_2_242<=Wgt_2_242; w_2_243<=Wgt_2_243; w_2_244<=Wgt_2_244; w_2_245<=Wgt_2_245; w_2_246<=Wgt_2_246; w_2_247<=Wgt_2_247; w_2_248<=Wgt_2_248; w_2_249<=Wgt_2_249; w_2_250<=Wgt_2_250; w_2_251<=Wgt_2_251; w_2_252<=Wgt_2_252; w_2_253<=Wgt_2_253; w_2_254<=Wgt_2_254; w_2_255<=Wgt_2_255; w_2_256<=Wgt_2_256; w_2_257<=Wgt_2_257; w_2_258<=Wgt_2_258; w_2_259<=Wgt_2_259; w_2_260<=Wgt_2_260; w_2_261<=Wgt_2_261; w_2_262<=Wgt_2_262; w_2_263<=Wgt_2_263; w_2_264<=Wgt_2_264; w_2_265<=Wgt_2_265; w_2_266<=Wgt_2_266; w_2_267<=Wgt_2_267; w_2_268<=Wgt_2_268; w_2_269<=Wgt_2_269; w_2_270<=Wgt_2_270; w_2_271<=Wgt_2_271; w_2_272<=Wgt_2_272; w_2_273<=Wgt_2_273; w_2_274<=Wgt_2_274; w_2_275<=Wgt_2_275; w_2_276<=Wgt_2_276; w_2_277<=Wgt_2_277; w_2_278<=Wgt_2_278; w_2_279<=Wgt_2_279; w_2_280<=Wgt_2_280; w_2_281<=Wgt_2_281; w_2_282<=Wgt_2_282; w_2_283<=Wgt_2_283; w_2_284<=Wgt_2_284; w_2_285<=Wgt_2_285; w_2_286<=Wgt_2_286; w_2_287<=Wgt_2_287; w_2_288<=Wgt_2_288; w_2_289<=Wgt_2_289; w_2_290<=Wgt_2_290; w_2_291<=Wgt_2_291; w_2_292<=Wgt_2_292; w_2_293<=Wgt_2_293; w_2_294<=Wgt_2_294; w_2_295<=Wgt_2_295; w_2_296<=Wgt_2_296; w_2_297<=Wgt_2_297; w_2_298<=Wgt_2_298; w_2_299<=Wgt_2_299; w_2_300<=Wgt_2_300; w_2_301<=Wgt_2_301; w_2_302<=Wgt_2_302; w_2_303<=Wgt_2_303; w_2_304<=Wgt_2_304; w_2_305<=Wgt_2_305; w_2_306<=Wgt_2_306; w_2_307<=Wgt_2_307; w_2_308<=Wgt_2_308; w_2_309<=Wgt_2_309; w_2_310<=Wgt_2_310; w_2_311<=Wgt_2_311; w_2_312<=Wgt_2_312; w_2_313<=Wgt_2_313; w_2_314<=Wgt_2_314; w_2_315<=Wgt_2_315; w_2_316<=Wgt_2_316; w_2_317<=Wgt_2_317; w_2_318<=Wgt_2_318; w_2_319<=Wgt_2_319; w_2_320<=Wgt_2_320; w_2_321<=Wgt_2_321; w_2_322<=Wgt_2_322; w_2_323<=Wgt_2_323; w_2_324<=Wgt_2_324; w_2_325<=Wgt_2_325; w_2_326<=Wgt_2_326; w_2_327<=Wgt_2_327; w_2_328<=Wgt_2_328; w_2_329<=Wgt_2_329; w_2_330<=Wgt_2_330; w_2_331<=Wgt_2_331; w_2_332<=Wgt_2_332; w_2_333<=Wgt_2_333; w_2_334<=Wgt_2_334; w_2_335<=Wgt_2_335; w_2_336<=Wgt_2_336; w_2_337<=Wgt_2_337; w_2_338<=Wgt_2_338; w_2_339<=Wgt_2_339; w_2_340<=Wgt_2_340; w_2_341<=Wgt_2_341; w_2_342<=Wgt_2_342; w_2_343<=Wgt_2_343; w_2_344<=Wgt_2_344; w_2_345<=Wgt_2_345; w_2_346<=Wgt_2_346; w_2_347<=Wgt_2_347; w_2_348<=Wgt_2_348; w_2_349<=Wgt_2_349; w_2_350<=Wgt_2_350; w_2_351<=Wgt_2_351; w_2_352<=Wgt_2_352; w_2_353<=Wgt_2_353; w_2_354<=Wgt_2_354; w_2_355<=Wgt_2_355; w_2_356<=Wgt_2_356; w_2_357<=Wgt_2_357; w_2_358<=Wgt_2_358; w_2_359<=Wgt_2_359; w_2_360<=Wgt_2_360; w_2_361<=Wgt_2_361; w_2_362<=Wgt_2_362; w_2_363<=Wgt_2_363; w_2_364<=Wgt_2_364; w_2_365<=Wgt_2_365; w_2_366<=Wgt_2_366; w_2_367<=Wgt_2_367; w_2_368<=Wgt_2_368; w_2_369<=Wgt_2_369; w_2_370<=Wgt_2_370; w_2_371<=Wgt_2_371; w_2_372<=Wgt_2_372; w_2_373<=Wgt_2_373; w_2_374<=Wgt_2_374; w_2_375<=Wgt_2_375; w_2_376<=Wgt_2_376; w_2_377<=Wgt_2_377; w_2_378<=Wgt_2_378; w_2_379<=Wgt_2_379; w_2_380<=Wgt_2_380; w_2_381<=Wgt_2_381; w_2_382<=Wgt_2_382; w_2_383<=Wgt_2_383; w_2_384<=Wgt_2_384; w_2_385<=Wgt_2_385; w_2_386<=Wgt_2_386; w_2_387<=Wgt_2_387; w_2_388<=Wgt_2_388; w_2_389<=Wgt_2_389; w_2_390<=Wgt_2_390; w_2_391<=Wgt_2_391; w_2_392<=Wgt_2_392; w_2_393<=Wgt_2_393; w_2_394<=Wgt_2_394; w_2_395<=Wgt_2_395; w_2_396<=Wgt_2_396; w_2_397<=Wgt_2_397; w_2_398<=Wgt_2_398; w_2_399<=Wgt_2_399; w_2_400<=Wgt_2_400; w_2_401<=Wgt_2_401; w_2_402<=Wgt_2_402; w_2_403<=Wgt_2_403; w_2_404<=Wgt_2_404; w_2_405<=Wgt_2_405; w_2_406<=Wgt_2_406; w_2_407<=Wgt_2_407; w_2_408<=Wgt_2_408; w_2_409<=Wgt_2_409; w_2_410<=Wgt_2_410; w_2_411<=Wgt_2_411; w_2_412<=Wgt_2_412; w_2_413<=Wgt_2_413; w_2_414<=Wgt_2_414; w_2_415<=Wgt_2_415; w_2_416<=Wgt_2_416; w_2_417<=Wgt_2_417; w_2_418<=Wgt_2_418; w_2_419<=Wgt_2_419; w_2_420<=Wgt_2_420; w_2_421<=Wgt_2_421; w_2_422<=Wgt_2_422; w_2_423<=Wgt_2_423; w_2_424<=Wgt_2_424; w_2_425<=Wgt_2_425; w_2_426<=Wgt_2_426; w_2_427<=Wgt_2_427; w_2_428<=Wgt_2_428; w_2_429<=Wgt_2_429; w_2_430<=Wgt_2_430; w_2_431<=Wgt_2_431; w_2_432<=Wgt_2_432; w_2_433<=Wgt_2_433; w_2_434<=Wgt_2_434; w_2_435<=Wgt_2_435; w_2_436<=Wgt_2_436; w_2_437<=Wgt_2_437; w_2_438<=Wgt_2_438; w_2_439<=Wgt_2_439; w_2_440<=Wgt_2_440; w_2_441<=Wgt_2_441; w_2_442<=Wgt_2_442; w_2_443<=Wgt_2_443; w_2_444<=Wgt_2_444; w_2_445<=Wgt_2_445; w_2_446<=Wgt_2_446; w_2_447<=Wgt_2_447; w_2_448<=Wgt_2_448; w_2_449<=Wgt_2_449; w_2_450<=Wgt_2_450; w_2_451<=Wgt_2_451; w_2_452<=Wgt_2_452; w_2_453<=Wgt_2_453; w_2_454<=Wgt_2_454; w_2_455<=Wgt_2_455; w_2_456<=Wgt_2_456; w_2_457<=Wgt_2_457; w_2_458<=Wgt_2_458; w_2_459<=Wgt_2_459; w_2_460<=Wgt_2_460; w_2_461<=Wgt_2_461; w_2_462<=Wgt_2_462; w_2_463<=Wgt_2_463; w_2_464<=Wgt_2_464; w_2_465<=Wgt_2_465; w_2_466<=Wgt_2_466; w_2_467<=Wgt_2_467; w_2_468<=Wgt_2_468; w_2_469<=Wgt_2_469; w_2_470<=Wgt_2_470; w_2_471<=Wgt_2_471; w_2_472<=Wgt_2_472; w_2_473<=Wgt_2_473; w_2_474<=Wgt_2_474; w_2_475<=Wgt_2_475; w_2_476<=Wgt_2_476; w_2_477<=Wgt_2_477; w_2_478<=Wgt_2_478; w_2_479<=Wgt_2_479; w_2_480<=Wgt_2_480; w_2_481<=Wgt_2_481; w_2_482<=Wgt_2_482; w_2_483<=Wgt_2_483; w_2_484<=Wgt_2_484; w_2_485<=Wgt_2_485; w_2_486<=Wgt_2_486; w_2_487<=Wgt_2_487; w_2_488<=Wgt_2_488; w_2_489<=Wgt_2_489; w_2_490<=Wgt_2_490; w_2_491<=Wgt_2_491; w_2_492<=Wgt_2_492; w_2_493<=Wgt_2_493; w_2_494<=Wgt_2_494; w_2_495<=Wgt_2_495; w_2_496<=Wgt_2_496; w_2_497<=Wgt_2_497; w_2_498<=Wgt_2_498; w_2_499<=Wgt_2_499; w_2_500<=Wgt_2_500; w_2_501<=Wgt_2_501; w_2_502<=Wgt_2_502; w_2_503<=Wgt_2_503; w_2_504<=Wgt_2_504; w_2_505<=Wgt_2_505; w_2_506<=Wgt_2_506; w_2_507<=Wgt_2_507; w_2_508<=Wgt_2_508; w_2_509<=Wgt_2_509; w_2_510<=Wgt_2_510; w_2_511<=Wgt_2_511; w_2_512<=Wgt_2_512; w_2_513<=Wgt_2_513; w_2_514<=Wgt_2_514; w_2_515<=Wgt_2_515; w_2_516<=Wgt_2_516; w_2_517<=Wgt_2_517; w_2_518<=Wgt_2_518; w_2_519<=Wgt_2_519; w_2_520<=Wgt_2_520; w_2_521<=Wgt_2_521; w_2_522<=Wgt_2_522; w_2_523<=Wgt_2_523; w_2_524<=Wgt_2_524; w_2_525<=Wgt_2_525; w_2_526<=Wgt_2_526; w_2_527<=Wgt_2_527; w_2_528<=Wgt_2_528; w_2_529<=Wgt_2_529; w_2_530<=Wgt_2_530; w_2_531<=Wgt_2_531; w_2_532<=Wgt_2_532; w_2_533<=Wgt_2_533; w_2_534<=Wgt_2_534; w_2_535<=Wgt_2_535; w_2_536<=Wgt_2_536; w_2_537<=Wgt_2_537; w_2_538<=Wgt_2_538; w_2_539<=Wgt_2_539; w_2_540<=Wgt_2_540; w_2_541<=Wgt_2_541; w_2_542<=Wgt_2_542; w_2_543<=Wgt_2_543; w_2_544<=Wgt_2_544; w_2_545<=Wgt_2_545; w_2_546<=Wgt_2_546; w_2_547<=Wgt_2_547; w_2_548<=Wgt_2_548; w_2_549<=Wgt_2_549; w_2_550<=Wgt_2_550; w_2_551<=Wgt_2_551; w_2_552<=Wgt_2_552; w_2_553<=Wgt_2_553; w_2_554<=Wgt_2_554; w_2_555<=Wgt_2_555; w_2_556<=Wgt_2_556; w_2_557<=Wgt_2_557; w_2_558<=Wgt_2_558; w_2_559<=Wgt_2_559; w_2_560<=Wgt_2_560; w_2_561<=Wgt_2_561; w_2_562<=Wgt_2_562; w_2_563<=Wgt_2_563; w_2_564<=Wgt_2_564; w_2_565<=Wgt_2_565; w_2_566<=Wgt_2_566; w_2_567<=Wgt_2_567; w_2_568<=Wgt_2_568; w_2_569<=Wgt_2_569; w_2_570<=Wgt_2_570; w_2_571<=Wgt_2_571; w_2_572<=Wgt_2_572; w_2_573<=Wgt_2_573; w_2_574<=Wgt_2_574; w_2_575<=Wgt_2_575; w_2_576<=Wgt_2_576; w_2_577<=Wgt_2_577; w_2_578<=Wgt_2_578; w_2_579<=Wgt_2_579; w_2_580<=Wgt_2_580; w_2_581<=Wgt_2_581; w_2_582<=Wgt_2_582; w_2_583<=Wgt_2_583; w_2_584<=Wgt_2_584; w_2_585<=Wgt_2_585; w_2_586<=Wgt_2_586; w_2_587<=Wgt_2_587; w_2_588<=Wgt_2_588; w_2_589<=Wgt_2_589; w_2_590<=Wgt_2_590; w_2_591<=Wgt_2_591; w_2_592<=Wgt_2_592; w_2_593<=Wgt_2_593; w_2_594<=Wgt_2_594; w_2_595<=Wgt_2_595; w_2_596<=Wgt_2_596; w_2_597<=Wgt_2_597; w_2_598<=Wgt_2_598; w_2_599<=Wgt_2_599; w_2_600<=Wgt_2_600; w_2_601<=Wgt_2_601; w_2_602<=Wgt_2_602; w_2_603<=Wgt_2_603; w_2_604<=Wgt_2_604; w_2_605<=Wgt_2_605; w_2_606<=Wgt_2_606; w_2_607<=Wgt_2_607; w_2_608<=Wgt_2_608; w_2_609<=Wgt_2_609; w_2_610<=Wgt_2_610; w_2_611<=Wgt_2_611; w_2_612<=Wgt_2_612; w_2_613<=Wgt_2_613; w_2_614<=Wgt_2_614; w_2_615<=Wgt_2_615; w_2_616<=Wgt_2_616; w_2_617<=Wgt_2_617; w_2_618<=Wgt_2_618; w_2_619<=Wgt_2_619; w_2_620<=Wgt_2_620; w_2_621<=Wgt_2_621; w_2_622<=Wgt_2_622; w_2_623<=Wgt_2_623; w_2_624<=Wgt_2_624; w_2_625<=Wgt_2_625; w_2_626<=Wgt_2_626; w_2_627<=Wgt_2_627; w_2_628<=Wgt_2_628; w_2_629<=Wgt_2_629; w_2_630<=Wgt_2_630; w_2_631<=Wgt_2_631; w_2_632<=Wgt_2_632; w_2_633<=Wgt_2_633; w_2_634<=Wgt_2_634; w_2_635<=Wgt_2_635; w_2_636<=Wgt_2_636; w_2_637<=Wgt_2_637; w_2_638<=Wgt_2_638; w_2_639<=Wgt_2_639; w_2_640<=Wgt_2_640; w_2_641<=Wgt_2_641; w_2_642<=Wgt_2_642; w_2_643<=Wgt_2_643; w_2_644<=Wgt_2_644; w_2_645<=Wgt_2_645; w_2_646<=Wgt_2_646; w_2_647<=Wgt_2_647; w_2_648<=Wgt_2_648; w_2_649<=Wgt_2_649; w_2_650<=Wgt_2_650; w_2_651<=Wgt_2_651; w_2_652<=Wgt_2_652; w_2_653<=Wgt_2_653; w_2_654<=Wgt_2_654; w_2_655<=Wgt_2_655; w_2_656<=Wgt_2_656; w_2_657<=Wgt_2_657; w_2_658<=Wgt_2_658; w_2_659<=Wgt_2_659; w_2_660<=Wgt_2_660; w_2_661<=Wgt_2_661; w_2_662<=Wgt_2_662; w_2_663<=Wgt_2_663; w_2_664<=Wgt_2_664; w_2_665<=Wgt_2_665; w_2_666<=Wgt_2_666; w_2_667<=Wgt_2_667; w_2_668<=Wgt_2_668; w_2_669<=Wgt_2_669; w_2_670<=Wgt_2_670; w_2_671<=Wgt_2_671; w_2_672<=Wgt_2_672; w_2_673<=Wgt_2_673; w_2_674<=Wgt_2_674; w_2_675<=Wgt_2_675; w_2_676<=Wgt_2_676; w_2_677<=Wgt_2_677; w_2_678<=Wgt_2_678; w_2_679<=Wgt_2_679; w_2_680<=Wgt_2_680; w_2_681<=Wgt_2_681; w_2_682<=Wgt_2_682; w_2_683<=Wgt_2_683; w_2_684<=Wgt_2_684; w_2_685<=Wgt_2_685; w_2_686<=Wgt_2_686; w_2_687<=Wgt_2_687; w_2_688<=Wgt_2_688; w_2_689<=Wgt_2_689; w_2_690<=Wgt_2_690; w_2_691<=Wgt_2_691; w_2_692<=Wgt_2_692; w_2_693<=Wgt_2_693; w_2_694<=Wgt_2_694; w_2_695<=Wgt_2_695; w_2_696<=Wgt_2_696; w_2_697<=Wgt_2_697; w_2_698<=Wgt_2_698; w_2_699<=Wgt_2_699; w_2_700<=Wgt_2_700; w_2_701<=Wgt_2_701; w_2_702<=Wgt_2_702; w_2_703<=Wgt_2_703; w_2_704<=Wgt_2_704; w_2_705<=Wgt_2_705; w_2_706<=Wgt_2_706; w_2_707<=Wgt_2_707; w_2_708<=Wgt_2_708; w_2_709<=Wgt_2_709; w_2_710<=Wgt_2_710; w_2_711<=Wgt_2_711; w_2_712<=Wgt_2_712; w_2_713<=Wgt_2_713; w_2_714<=Wgt_2_714; w_2_715<=Wgt_2_715; w_2_716<=Wgt_2_716; w_2_717<=Wgt_2_717; w_2_718<=Wgt_2_718; w_2_719<=Wgt_2_719; w_2_720<=Wgt_2_720; w_2_721<=Wgt_2_721; w_2_722<=Wgt_2_722; w_2_723<=Wgt_2_723; w_2_724<=Wgt_2_724; w_2_725<=Wgt_2_725; w_2_726<=Wgt_2_726; w_2_727<=Wgt_2_727; w_2_728<=Wgt_2_728; w_2_729<=Wgt_2_729; w_2_730<=Wgt_2_730; w_2_731<=Wgt_2_731; w_2_732<=Wgt_2_732; w_2_733<=Wgt_2_733; w_2_734<=Wgt_2_734; w_2_735<=Wgt_2_735; w_2_736<=Wgt_2_736; w_2_737<=Wgt_2_737; w_2_738<=Wgt_2_738; w_2_739<=Wgt_2_739; w_2_740<=Wgt_2_740; w_2_741<=Wgt_2_741; w_2_742<=Wgt_2_742; w_2_743<=Wgt_2_743; w_2_744<=Wgt_2_744; w_2_745<=Wgt_2_745; w_2_746<=Wgt_2_746; w_2_747<=Wgt_2_747; w_2_748<=Wgt_2_748; w_2_749<=Wgt_2_749; w_2_750<=Wgt_2_750; w_2_751<=Wgt_2_751; w_2_752<=Wgt_2_752; w_2_753<=Wgt_2_753; w_2_754<=Wgt_2_754; w_2_755<=Wgt_2_755; w_2_756<=Wgt_2_756; w_2_757<=Wgt_2_757; w_2_758<=Wgt_2_758; w_2_759<=Wgt_2_759; w_2_760<=Wgt_2_760; w_2_761<=Wgt_2_761; w_2_762<=Wgt_2_762; w_2_763<=Wgt_2_763; w_2_764<=Wgt_2_764; w_2_765<=Wgt_2_765; w_2_766<=Wgt_2_766; w_2_767<=Wgt_2_767; w_2_768<=Wgt_2_768; w_2_769<=Wgt_2_769; w_2_770<=Wgt_2_770; w_2_771<=Wgt_2_771; w_2_772<=Wgt_2_772; w_2_773<=Wgt_2_773; w_2_774<=Wgt_2_774; w_2_775<=Wgt_2_775; w_2_776<=Wgt_2_776; w_2_777<=Wgt_2_777; w_2_778<=Wgt_2_778; w_2_779<=Wgt_2_779; w_2_780<=Wgt_2_780; w_2_781<=Wgt_2_781; w_2_782<=Wgt_2_782; w_2_783<=Wgt_2_783; w_2_784<=Wgt_2_784; 
					w_3_0<=Wgt_3_0; w_3_1<=Wgt_3_1; w_3_2<=Wgt_3_2; w_3_3<=Wgt_3_3; w_3_4<=Wgt_3_4; w_3_5<=Wgt_3_5; w_3_6<=Wgt_3_6; w_3_7<=Wgt_3_7; w_3_8<=Wgt_3_8; w_3_9<=Wgt_3_9; w_3_10<=Wgt_3_10; w_3_11<=Wgt_3_11; w_3_12<=Wgt_3_12; w_3_13<=Wgt_3_13; w_3_14<=Wgt_3_14; w_3_15<=Wgt_3_15; w_3_16<=Wgt_3_16; w_3_17<=Wgt_3_17; w_3_18<=Wgt_3_18; w_3_19<=Wgt_3_19; w_3_20<=Wgt_3_20; w_3_21<=Wgt_3_21; w_3_22<=Wgt_3_22; w_3_23<=Wgt_3_23; w_3_24<=Wgt_3_24; w_3_25<=Wgt_3_25; w_3_26<=Wgt_3_26; w_3_27<=Wgt_3_27; w_3_28<=Wgt_3_28; w_3_29<=Wgt_3_29; w_3_30<=Wgt_3_30; w_3_31<=Wgt_3_31; w_3_32<=Wgt_3_32; w_3_33<=Wgt_3_33; w_3_34<=Wgt_3_34; w_3_35<=Wgt_3_35; w_3_36<=Wgt_3_36; w_3_37<=Wgt_3_37; w_3_38<=Wgt_3_38; w_3_39<=Wgt_3_39; w_3_40<=Wgt_3_40; w_3_41<=Wgt_3_41; w_3_42<=Wgt_3_42; w_3_43<=Wgt_3_43; w_3_44<=Wgt_3_44; w_3_45<=Wgt_3_45; w_3_46<=Wgt_3_46; w_3_47<=Wgt_3_47; w_3_48<=Wgt_3_48; w_3_49<=Wgt_3_49; w_3_50<=Wgt_3_50; w_3_51<=Wgt_3_51; w_3_52<=Wgt_3_52; w_3_53<=Wgt_3_53; w_3_54<=Wgt_3_54; w_3_55<=Wgt_3_55; w_3_56<=Wgt_3_56; w_3_57<=Wgt_3_57; w_3_58<=Wgt_3_58; w_3_59<=Wgt_3_59; w_3_60<=Wgt_3_60; w_3_61<=Wgt_3_61; w_3_62<=Wgt_3_62; w_3_63<=Wgt_3_63; w_3_64<=Wgt_3_64; w_3_65<=Wgt_3_65; w_3_66<=Wgt_3_66; w_3_67<=Wgt_3_67; w_3_68<=Wgt_3_68; w_3_69<=Wgt_3_69; w_3_70<=Wgt_3_70; w_3_71<=Wgt_3_71; w_3_72<=Wgt_3_72; w_3_73<=Wgt_3_73; w_3_74<=Wgt_3_74; w_3_75<=Wgt_3_75; w_3_76<=Wgt_3_76; w_3_77<=Wgt_3_77; w_3_78<=Wgt_3_78; w_3_79<=Wgt_3_79; w_3_80<=Wgt_3_80; w_3_81<=Wgt_3_81; w_3_82<=Wgt_3_82; w_3_83<=Wgt_3_83; w_3_84<=Wgt_3_84; w_3_85<=Wgt_3_85; w_3_86<=Wgt_3_86; w_3_87<=Wgt_3_87; w_3_88<=Wgt_3_88; w_3_89<=Wgt_3_89; w_3_90<=Wgt_3_90; w_3_91<=Wgt_3_91; w_3_92<=Wgt_3_92; w_3_93<=Wgt_3_93; w_3_94<=Wgt_3_94; w_3_95<=Wgt_3_95; w_3_96<=Wgt_3_96; w_3_97<=Wgt_3_97; w_3_98<=Wgt_3_98; w_3_99<=Wgt_3_99; w_3_100<=Wgt_3_100; w_3_101<=Wgt_3_101; w_3_102<=Wgt_3_102; w_3_103<=Wgt_3_103; w_3_104<=Wgt_3_104; w_3_105<=Wgt_3_105; w_3_106<=Wgt_3_106; w_3_107<=Wgt_3_107; w_3_108<=Wgt_3_108; w_3_109<=Wgt_3_109; w_3_110<=Wgt_3_110; w_3_111<=Wgt_3_111; w_3_112<=Wgt_3_112; w_3_113<=Wgt_3_113; w_3_114<=Wgt_3_114; w_3_115<=Wgt_3_115; w_3_116<=Wgt_3_116; w_3_117<=Wgt_3_117; w_3_118<=Wgt_3_118; w_3_119<=Wgt_3_119; w_3_120<=Wgt_3_120; w_3_121<=Wgt_3_121; w_3_122<=Wgt_3_122; w_3_123<=Wgt_3_123; w_3_124<=Wgt_3_124; w_3_125<=Wgt_3_125; w_3_126<=Wgt_3_126; w_3_127<=Wgt_3_127; w_3_128<=Wgt_3_128; w_3_129<=Wgt_3_129; w_3_130<=Wgt_3_130; w_3_131<=Wgt_3_131; w_3_132<=Wgt_3_132; w_3_133<=Wgt_3_133; w_3_134<=Wgt_3_134; w_3_135<=Wgt_3_135; w_3_136<=Wgt_3_136; w_3_137<=Wgt_3_137; w_3_138<=Wgt_3_138; w_3_139<=Wgt_3_139; w_3_140<=Wgt_3_140; w_3_141<=Wgt_3_141; w_3_142<=Wgt_3_142; w_3_143<=Wgt_3_143; w_3_144<=Wgt_3_144; w_3_145<=Wgt_3_145; w_3_146<=Wgt_3_146; w_3_147<=Wgt_3_147; w_3_148<=Wgt_3_148; w_3_149<=Wgt_3_149; w_3_150<=Wgt_3_150; w_3_151<=Wgt_3_151; w_3_152<=Wgt_3_152; w_3_153<=Wgt_3_153; w_3_154<=Wgt_3_154; w_3_155<=Wgt_3_155; w_3_156<=Wgt_3_156; w_3_157<=Wgt_3_157; w_3_158<=Wgt_3_158; w_3_159<=Wgt_3_159; w_3_160<=Wgt_3_160; w_3_161<=Wgt_3_161; w_3_162<=Wgt_3_162; w_3_163<=Wgt_3_163; w_3_164<=Wgt_3_164; w_3_165<=Wgt_3_165; w_3_166<=Wgt_3_166; w_3_167<=Wgt_3_167; w_3_168<=Wgt_3_168; w_3_169<=Wgt_3_169; w_3_170<=Wgt_3_170; w_3_171<=Wgt_3_171; w_3_172<=Wgt_3_172; w_3_173<=Wgt_3_173; w_3_174<=Wgt_3_174; w_3_175<=Wgt_3_175; w_3_176<=Wgt_3_176; w_3_177<=Wgt_3_177; w_3_178<=Wgt_3_178; w_3_179<=Wgt_3_179; w_3_180<=Wgt_3_180; w_3_181<=Wgt_3_181; w_3_182<=Wgt_3_182; w_3_183<=Wgt_3_183; w_3_184<=Wgt_3_184; w_3_185<=Wgt_3_185; w_3_186<=Wgt_3_186; w_3_187<=Wgt_3_187; w_3_188<=Wgt_3_188; w_3_189<=Wgt_3_189; w_3_190<=Wgt_3_190; w_3_191<=Wgt_3_191; w_3_192<=Wgt_3_192; w_3_193<=Wgt_3_193; w_3_194<=Wgt_3_194; w_3_195<=Wgt_3_195; w_3_196<=Wgt_3_196; w_3_197<=Wgt_3_197; w_3_198<=Wgt_3_198; w_3_199<=Wgt_3_199; w_3_200<=Wgt_3_200; w_3_201<=Wgt_3_201; w_3_202<=Wgt_3_202; w_3_203<=Wgt_3_203; w_3_204<=Wgt_3_204; w_3_205<=Wgt_3_205; w_3_206<=Wgt_3_206; w_3_207<=Wgt_3_207; w_3_208<=Wgt_3_208; w_3_209<=Wgt_3_209; w_3_210<=Wgt_3_210; w_3_211<=Wgt_3_211; w_3_212<=Wgt_3_212; w_3_213<=Wgt_3_213; w_3_214<=Wgt_3_214; w_3_215<=Wgt_3_215; w_3_216<=Wgt_3_216; w_3_217<=Wgt_3_217; w_3_218<=Wgt_3_218; w_3_219<=Wgt_3_219; w_3_220<=Wgt_3_220; w_3_221<=Wgt_3_221; w_3_222<=Wgt_3_222; w_3_223<=Wgt_3_223; w_3_224<=Wgt_3_224; w_3_225<=Wgt_3_225; w_3_226<=Wgt_3_226; w_3_227<=Wgt_3_227; w_3_228<=Wgt_3_228; w_3_229<=Wgt_3_229; w_3_230<=Wgt_3_230; w_3_231<=Wgt_3_231; w_3_232<=Wgt_3_232; w_3_233<=Wgt_3_233; w_3_234<=Wgt_3_234; w_3_235<=Wgt_3_235; w_3_236<=Wgt_3_236; w_3_237<=Wgt_3_237; w_3_238<=Wgt_3_238; w_3_239<=Wgt_3_239; w_3_240<=Wgt_3_240; w_3_241<=Wgt_3_241; w_3_242<=Wgt_3_242; w_3_243<=Wgt_3_243; w_3_244<=Wgt_3_244; w_3_245<=Wgt_3_245; w_3_246<=Wgt_3_246; w_3_247<=Wgt_3_247; w_3_248<=Wgt_3_248; w_3_249<=Wgt_3_249; w_3_250<=Wgt_3_250; w_3_251<=Wgt_3_251; w_3_252<=Wgt_3_252; w_3_253<=Wgt_3_253; w_3_254<=Wgt_3_254; w_3_255<=Wgt_3_255; w_3_256<=Wgt_3_256; w_3_257<=Wgt_3_257; w_3_258<=Wgt_3_258; w_3_259<=Wgt_3_259; w_3_260<=Wgt_3_260; w_3_261<=Wgt_3_261; w_3_262<=Wgt_3_262; w_3_263<=Wgt_3_263; w_3_264<=Wgt_3_264; w_3_265<=Wgt_3_265; w_3_266<=Wgt_3_266; w_3_267<=Wgt_3_267; w_3_268<=Wgt_3_268; w_3_269<=Wgt_3_269; w_3_270<=Wgt_3_270; w_3_271<=Wgt_3_271; w_3_272<=Wgt_3_272; w_3_273<=Wgt_3_273; w_3_274<=Wgt_3_274; w_3_275<=Wgt_3_275; w_3_276<=Wgt_3_276; w_3_277<=Wgt_3_277; w_3_278<=Wgt_3_278; w_3_279<=Wgt_3_279; w_3_280<=Wgt_3_280; w_3_281<=Wgt_3_281; w_3_282<=Wgt_3_282; w_3_283<=Wgt_3_283; w_3_284<=Wgt_3_284; w_3_285<=Wgt_3_285; w_3_286<=Wgt_3_286; w_3_287<=Wgt_3_287; w_3_288<=Wgt_3_288; w_3_289<=Wgt_3_289; w_3_290<=Wgt_3_290; w_3_291<=Wgt_3_291; w_3_292<=Wgt_3_292; w_3_293<=Wgt_3_293; w_3_294<=Wgt_3_294; w_3_295<=Wgt_3_295; w_3_296<=Wgt_3_296; w_3_297<=Wgt_3_297; w_3_298<=Wgt_3_298; w_3_299<=Wgt_3_299; w_3_300<=Wgt_3_300; w_3_301<=Wgt_3_301; w_3_302<=Wgt_3_302; w_3_303<=Wgt_3_303; w_3_304<=Wgt_3_304; w_3_305<=Wgt_3_305; w_3_306<=Wgt_3_306; w_3_307<=Wgt_3_307; w_3_308<=Wgt_3_308; w_3_309<=Wgt_3_309; w_3_310<=Wgt_3_310; w_3_311<=Wgt_3_311; w_3_312<=Wgt_3_312; w_3_313<=Wgt_3_313; w_3_314<=Wgt_3_314; w_3_315<=Wgt_3_315; w_3_316<=Wgt_3_316; w_3_317<=Wgt_3_317; w_3_318<=Wgt_3_318; w_3_319<=Wgt_3_319; w_3_320<=Wgt_3_320; w_3_321<=Wgt_3_321; w_3_322<=Wgt_3_322; w_3_323<=Wgt_3_323; w_3_324<=Wgt_3_324; w_3_325<=Wgt_3_325; w_3_326<=Wgt_3_326; w_3_327<=Wgt_3_327; w_3_328<=Wgt_3_328; w_3_329<=Wgt_3_329; w_3_330<=Wgt_3_330; w_3_331<=Wgt_3_331; w_3_332<=Wgt_3_332; w_3_333<=Wgt_3_333; w_3_334<=Wgt_3_334; w_3_335<=Wgt_3_335; w_3_336<=Wgt_3_336; w_3_337<=Wgt_3_337; w_3_338<=Wgt_3_338; w_3_339<=Wgt_3_339; w_3_340<=Wgt_3_340; w_3_341<=Wgt_3_341; w_3_342<=Wgt_3_342; w_3_343<=Wgt_3_343; w_3_344<=Wgt_3_344; w_3_345<=Wgt_3_345; w_3_346<=Wgt_3_346; w_3_347<=Wgt_3_347; w_3_348<=Wgt_3_348; w_3_349<=Wgt_3_349; w_3_350<=Wgt_3_350; w_3_351<=Wgt_3_351; w_3_352<=Wgt_3_352; w_3_353<=Wgt_3_353; w_3_354<=Wgt_3_354; w_3_355<=Wgt_3_355; w_3_356<=Wgt_3_356; w_3_357<=Wgt_3_357; w_3_358<=Wgt_3_358; w_3_359<=Wgt_3_359; w_3_360<=Wgt_3_360; w_3_361<=Wgt_3_361; w_3_362<=Wgt_3_362; w_3_363<=Wgt_3_363; w_3_364<=Wgt_3_364; w_3_365<=Wgt_3_365; w_3_366<=Wgt_3_366; w_3_367<=Wgt_3_367; w_3_368<=Wgt_3_368; w_3_369<=Wgt_3_369; w_3_370<=Wgt_3_370; w_3_371<=Wgt_3_371; w_3_372<=Wgt_3_372; w_3_373<=Wgt_3_373; w_3_374<=Wgt_3_374; w_3_375<=Wgt_3_375; w_3_376<=Wgt_3_376; w_3_377<=Wgt_3_377; w_3_378<=Wgt_3_378; w_3_379<=Wgt_3_379; w_3_380<=Wgt_3_380; w_3_381<=Wgt_3_381; w_3_382<=Wgt_3_382; w_3_383<=Wgt_3_383; w_3_384<=Wgt_3_384; w_3_385<=Wgt_3_385; w_3_386<=Wgt_3_386; w_3_387<=Wgt_3_387; w_3_388<=Wgt_3_388; w_3_389<=Wgt_3_389; w_3_390<=Wgt_3_390; w_3_391<=Wgt_3_391; w_3_392<=Wgt_3_392; w_3_393<=Wgt_3_393; w_3_394<=Wgt_3_394; w_3_395<=Wgt_3_395; w_3_396<=Wgt_3_396; w_3_397<=Wgt_3_397; w_3_398<=Wgt_3_398; w_3_399<=Wgt_3_399; w_3_400<=Wgt_3_400; w_3_401<=Wgt_3_401; w_3_402<=Wgt_3_402; w_3_403<=Wgt_3_403; w_3_404<=Wgt_3_404; w_3_405<=Wgt_3_405; w_3_406<=Wgt_3_406; w_3_407<=Wgt_3_407; w_3_408<=Wgt_3_408; w_3_409<=Wgt_3_409; w_3_410<=Wgt_3_410; w_3_411<=Wgt_3_411; w_3_412<=Wgt_3_412; w_3_413<=Wgt_3_413; w_3_414<=Wgt_3_414; w_3_415<=Wgt_3_415; w_3_416<=Wgt_3_416; w_3_417<=Wgt_3_417; w_3_418<=Wgt_3_418; w_3_419<=Wgt_3_419; w_3_420<=Wgt_3_420; w_3_421<=Wgt_3_421; w_3_422<=Wgt_3_422; w_3_423<=Wgt_3_423; w_3_424<=Wgt_3_424; w_3_425<=Wgt_3_425; w_3_426<=Wgt_3_426; w_3_427<=Wgt_3_427; w_3_428<=Wgt_3_428; w_3_429<=Wgt_3_429; w_3_430<=Wgt_3_430; w_3_431<=Wgt_3_431; w_3_432<=Wgt_3_432; w_3_433<=Wgt_3_433; w_3_434<=Wgt_3_434; w_3_435<=Wgt_3_435; w_3_436<=Wgt_3_436; w_3_437<=Wgt_3_437; w_3_438<=Wgt_3_438; w_3_439<=Wgt_3_439; w_3_440<=Wgt_3_440; w_3_441<=Wgt_3_441; w_3_442<=Wgt_3_442; w_3_443<=Wgt_3_443; w_3_444<=Wgt_3_444; w_3_445<=Wgt_3_445; w_3_446<=Wgt_3_446; w_3_447<=Wgt_3_447; w_3_448<=Wgt_3_448; w_3_449<=Wgt_3_449; w_3_450<=Wgt_3_450; w_3_451<=Wgt_3_451; w_3_452<=Wgt_3_452; w_3_453<=Wgt_3_453; w_3_454<=Wgt_3_454; w_3_455<=Wgt_3_455; w_3_456<=Wgt_3_456; w_3_457<=Wgt_3_457; w_3_458<=Wgt_3_458; w_3_459<=Wgt_3_459; w_3_460<=Wgt_3_460; w_3_461<=Wgt_3_461; w_3_462<=Wgt_3_462; w_3_463<=Wgt_3_463; w_3_464<=Wgt_3_464; w_3_465<=Wgt_3_465; w_3_466<=Wgt_3_466; w_3_467<=Wgt_3_467; w_3_468<=Wgt_3_468; w_3_469<=Wgt_3_469; w_3_470<=Wgt_3_470; w_3_471<=Wgt_3_471; w_3_472<=Wgt_3_472; w_3_473<=Wgt_3_473; w_3_474<=Wgt_3_474; w_3_475<=Wgt_3_475; w_3_476<=Wgt_3_476; w_3_477<=Wgt_3_477; w_3_478<=Wgt_3_478; w_3_479<=Wgt_3_479; w_3_480<=Wgt_3_480; w_3_481<=Wgt_3_481; w_3_482<=Wgt_3_482; w_3_483<=Wgt_3_483; w_3_484<=Wgt_3_484; w_3_485<=Wgt_3_485; w_3_486<=Wgt_3_486; w_3_487<=Wgt_3_487; w_3_488<=Wgt_3_488; w_3_489<=Wgt_3_489; w_3_490<=Wgt_3_490; w_3_491<=Wgt_3_491; w_3_492<=Wgt_3_492; w_3_493<=Wgt_3_493; w_3_494<=Wgt_3_494; w_3_495<=Wgt_3_495; w_3_496<=Wgt_3_496; w_3_497<=Wgt_3_497; w_3_498<=Wgt_3_498; w_3_499<=Wgt_3_499; w_3_500<=Wgt_3_500; w_3_501<=Wgt_3_501; w_3_502<=Wgt_3_502; w_3_503<=Wgt_3_503; w_3_504<=Wgt_3_504; w_3_505<=Wgt_3_505; w_3_506<=Wgt_3_506; w_3_507<=Wgt_3_507; w_3_508<=Wgt_3_508; w_3_509<=Wgt_3_509; w_3_510<=Wgt_3_510; w_3_511<=Wgt_3_511; w_3_512<=Wgt_3_512; w_3_513<=Wgt_3_513; w_3_514<=Wgt_3_514; w_3_515<=Wgt_3_515; w_3_516<=Wgt_3_516; w_3_517<=Wgt_3_517; w_3_518<=Wgt_3_518; w_3_519<=Wgt_3_519; w_3_520<=Wgt_3_520; w_3_521<=Wgt_3_521; w_3_522<=Wgt_3_522; w_3_523<=Wgt_3_523; w_3_524<=Wgt_3_524; w_3_525<=Wgt_3_525; w_3_526<=Wgt_3_526; w_3_527<=Wgt_3_527; w_3_528<=Wgt_3_528; w_3_529<=Wgt_3_529; w_3_530<=Wgt_3_530; w_3_531<=Wgt_3_531; w_3_532<=Wgt_3_532; w_3_533<=Wgt_3_533; w_3_534<=Wgt_3_534; w_3_535<=Wgt_3_535; w_3_536<=Wgt_3_536; w_3_537<=Wgt_3_537; w_3_538<=Wgt_3_538; w_3_539<=Wgt_3_539; w_3_540<=Wgt_3_540; w_3_541<=Wgt_3_541; w_3_542<=Wgt_3_542; w_3_543<=Wgt_3_543; w_3_544<=Wgt_3_544; w_3_545<=Wgt_3_545; w_3_546<=Wgt_3_546; w_3_547<=Wgt_3_547; w_3_548<=Wgt_3_548; w_3_549<=Wgt_3_549; w_3_550<=Wgt_3_550; w_3_551<=Wgt_3_551; w_3_552<=Wgt_3_552; w_3_553<=Wgt_3_553; w_3_554<=Wgt_3_554; w_3_555<=Wgt_3_555; w_3_556<=Wgt_3_556; w_3_557<=Wgt_3_557; w_3_558<=Wgt_3_558; w_3_559<=Wgt_3_559; w_3_560<=Wgt_3_560; w_3_561<=Wgt_3_561; w_3_562<=Wgt_3_562; w_3_563<=Wgt_3_563; w_3_564<=Wgt_3_564; w_3_565<=Wgt_3_565; w_3_566<=Wgt_3_566; w_3_567<=Wgt_3_567; w_3_568<=Wgt_3_568; w_3_569<=Wgt_3_569; w_3_570<=Wgt_3_570; w_3_571<=Wgt_3_571; w_3_572<=Wgt_3_572; w_3_573<=Wgt_3_573; w_3_574<=Wgt_3_574; w_3_575<=Wgt_3_575; w_3_576<=Wgt_3_576; w_3_577<=Wgt_3_577; w_3_578<=Wgt_3_578; w_3_579<=Wgt_3_579; w_3_580<=Wgt_3_580; w_3_581<=Wgt_3_581; w_3_582<=Wgt_3_582; w_3_583<=Wgt_3_583; w_3_584<=Wgt_3_584; w_3_585<=Wgt_3_585; w_3_586<=Wgt_3_586; w_3_587<=Wgt_3_587; w_3_588<=Wgt_3_588; w_3_589<=Wgt_3_589; w_3_590<=Wgt_3_590; w_3_591<=Wgt_3_591; w_3_592<=Wgt_3_592; w_3_593<=Wgt_3_593; w_3_594<=Wgt_3_594; w_3_595<=Wgt_3_595; w_3_596<=Wgt_3_596; w_3_597<=Wgt_3_597; w_3_598<=Wgt_3_598; w_3_599<=Wgt_3_599; w_3_600<=Wgt_3_600; w_3_601<=Wgt_3_601; w_3_602<=Wgt_3_602; w_3_603<=Wgt_3_603; w_3_604<=Wgt_3_604; w_3_605<=Wgt_3_605; w_3_606<=Wgt_3_606; w_3_607<=Wgt_3_607; w_3_608<=Wgt_3_608; w_3_609<=Wgt_3_609; w_3_610<=Wgt_3_610; w_3_611<=Wgt_3_611; w_3_612<=Wgt_3_612; w_3_613<=Wgt_3_613; w_3_614<=Wgt_3_614; w_3_615<=Wgt_3_615; w_3_616<=Wgt_3_616; w_3_617<=Wgt_3_617; w_3_618<=Wgt_3_618; w_3_619<=Wgt_3_619; w_3_620<=Wgt_3_620; w_3_621<=Wgt_3_621; w_3_622<=Wgt_3_622; w_3_623<=Wgt_3_623; w_3_624<=Wgt_3_624; w_3_625<=Wgt_3_625; w_3_626<=Wgt_3_626; w_3_627<=Wgt_3_627; w_3_628<=Wgt_3_628; w_3_629<=Wgt_3_629; w_3_630<=Wgt_3_630; w_3_631<=Wgt_3_631; w_3_632<=Wgt_3_632; w_3_633<=Wgt_3_633; w_3_634<=Wgt_3_634; w_3_635<=Wgt_3_635; w_3_636<=Wgt_3_636; w_3_637<=Wgt_3_637; w_3_638<=Wgt_3_638; w_3_639<=Wgt_3_639; w_3_640<=Wgt_3_640; w_3_641<=Wgt_3_641; w_3_642<=Wgt_3_642; w_3_643<=Wgt_3_643; w_3_644<=Wgt_3_644; w_3_645<=Wgt_3_645; w_3_646<=Wgt_3_646; w_3_647<=Wgt_3_647; w_3_648<=Wgt_3_648; w_3_649<=Wgt_3_649; w_3_650<=Wgt_3_650; w_3_651<=Wgt_3_651; w_3_652<=Wgt_3_652; w_3_653<=Wgt_3_653; w_3_654<=Wgt_3_654; w_3_655<=Wgt_3_655; w_3_656<=Wgt_3_656; w_3_657<=Wgt_3_657; w_3_658<=Wgt_3_658; w_3_659<=Wgt_3_659; w_3_660<=Wgt_3_660; w_3_661<=Wgt_3_661; w_3_662<=Wgt_3_662; w_3_663<=Wgt_3_663; w_3_664<=Wgt_3_664; w_3_665<=Wgt_3_665; w_3_666<=Wgt_3_666; w_3_667<=Wgt_3_667; w_3_668<=Wgt_3_668; w_3_669<=Wgt_3_669; w_3_670<=Wgt_3_670; w_3_671<=Wgt_3_671; w_3_672<=Wgt_3_672; w_3_673<=Wgt_3_673; w_3_674<=Wgt_3_674; w_3_675<=Wgt_3_675; w_3_676<=Wgt_3_676; w_3_677<=Wgt_3_677; w_3_678<=Wgt_3_678; w_3_679<=Wgt_3_679; w_3_680<=Wgt_3_680; w_3_681<=Wgt_3_681; w_3_682<=Wgt_3_682; w_3_683<=Wgt_3_683; w_3_684<=Wgt_3_684; w_3_685<=Wgt_3_685; w_3_686<=Wgt_3_686; w_3_687<=Wgt_3_687; w_3_688<=Wgt_3_688; w_3_689<=Wgt_3_689; w_3_690<=Wgt_3_690; w_3_691<=Wgt_3_691; w_3_692<=Wgt_3_692; w_3_693<=Wgt_3_693; w_3_694<=Wgt_3_694; w_3_695<=Wgt_3_695; w_3_696<=Wgt_3_696; w_3_697<=Wgt_3_697; w_3_698<=Wgt_3_698; w_3_699<=Wgt_3_699; w_3_700<=Wgt_3_700; w_3_701<=Wgt_3_701; w_3_702<=Wgt_3_702; w_3_703<=Wgt_3_703; w_3_704<=Wgt_3_704; w_3_705<=Wgt_3_705; w_3_706<=Wgt_3_706; w_3_707<=Wgt_3_707; w_3_708<=Wgt_3_708; w_3_709<=Wgt_3_709; w_3_710<=Wgt_3_710; w_3_711<=Wgt_3_711; w_3_712<=Wgt_3_712; w_3_713<=Wgt_3_713; w_3_714<=Wgt_3_714; w_3_715<=Wgt_3_715; w_3_716<=Wgt_3_716; w_3_717<=Wgt_3_717; w_3_718<=Wgt_3_718; w_3_719<=Wgt_3_719; w_3_720<=Wgt_3_720; w_3_721<=Wgt_3_721; w_3_722<=Wgt_3_722; w_3_723<=Wgt_3_723; w_3_724<=Wgt_3_724; w_3_725<=Wgt_3_725; w_3_726<=Wgt_3_726; w_3_727<=Wgt_3_727; w_3_728<=Wgt_3_728; w_3_729<=Wgt_3_729; w_3_730<=Wgt_3_730; w_3_731<=Wgt_3_731; w_3_732<=Wgt_3_732; w_3_733<=Wgt_3_733; w_3_734<=Wgt_3_734; w_3_735<=Wgt_3_735; w_3_736<=Wgt_3_736; w_3_737<=Wgt_3_737; w_3_738<=Wgt_3_738; w_3_739<=Wgt_3_739; w_3_740<=Wgt_3_740; w_3_741<=Wgt_3_741; w_3_742<=Wgt_3_742; w_3_743<=Wgt_3_743; w_3_744<=Wgt_3_744; w_3_745<=Wgt_3_745; w_3_746<=Wgt_3_746; w_3_747<=Wgt_3_747; w_3_748<=Wgt_3_748; w_3_749<=Wgt_3_749; w_3_750<=Wgt_3_750; w_3_751<=Wgt_3_751; w_3_752<=Wgt_3_752; w_3_753<=Wgt_3_753; w_3_754<=Wgt_3_754; w_3_755<=Wgt_3_755; w_3_756<=Wgt_3_756; w_3_757<=Wgt_3_757; w_3_758<=Wgt_3_758; w_3_759<=Wgt_3_759; w_3_760<=Wgt_3_760; w_3_761<=Wgt_3_761; w_3_762<=Wgt_3_762; w_3_763<=Wgt_3_763; w_3_764<=Wgt_3_764; w_3_765<=Wgt_3_765; w_3_766<=Wgt_3_766; w_3_767<=Wgt_3_767; w_3_768<=Wgt_3_768; w_3_769<=Wgt_3_769; w_3_770<=Wgt_3_770; w_3_771<=Wgt_3_771; w_3_772<=Wgt_3_772; w_3_773<=Wgt_3_773; w_3_774<=Wgt_3_774; w_3_775<=Wgt_3_775; w_3_776<=Wgt_3_776; w_3_777<=Wgt_3_777; w_3_778<=Wgt_3_778; w_3_779<=Wgt_3_779; w_3_780<=Wgt_3_780; w_3_781<=Wgt_3_781; w_3_782<=Wgt_3_782; w_3_783<=Wgt_3_783; w_3_784<=Wgt_3_784; 
					w_4_0<=Wgt_4_0; w_4_1<=Wgt_4_1; w_4_2<=Wgt_4_2; w_4_3<=Wgt_4_3; w_4_4<=Wgt_4_4; w_4_5<=Wgt_4_5; w_4_6<=Wgt_4_6; w_4_7<=Wgt_4_7; w_4_8<=Wgt_4_8; w_4_9<=Wgt_4_9; w_4_10<=Wgt_4_10; w_4_11<=Wgt_4_11; w_4_12<=Wgt_4_12; w_4_13<=Wgt_4_13; w_4_14<=Wgt_4_14; w_4_15<=Wgt_4_15; w_4_16<=Wgt_4_16; w_4_17<=Wgt_4_17; w_4_18<=Wgt_4_18; w_4_19<=Wgt_4_19; w_4_20<=Wgt_4_20; w_4_21<=Wgt_4_21; w_4_22<=Wgt_4_22; w_4_23<=Wgt_4_23; w_4_24<=Wgt_4_24; w_4_25<=Wgt_4_25; w_4_26<=Wgt_4_26; w_4_27<=Wgt_4_27; w_4_28<=Wgt_4_28; w_4_29<=Wgt_4_29; w_4_30<=Wgt_4_30; w_4_31<=Wgt_4_31; w_4_32<=Wgt_4_32; w_4_33<=Wgt_4_33; w_4_34<=Wgt_4_34; w_4_35<=Wgt_4_35; w_4_36<=Wgt_4_36; w_4_37<=Wgt_4_37; w_4_38<=Wgt_4_38; w_4_39<=Wgt_4_39; w_4_40<=Wgt_4_40; w_4_41<=Wgt_4_41; w_4_42<=Wgt_4_42; w_4_43<=Wgt_4_43; w_4_44<=Wgt_4_44; w_4_45<=Wgt_4_45; w_4_46<=Wgt_4_46; w_4_47<=Wgt_4_47; w_4_48<=Wgt_4_48; w_4_49<=Wgt_4_49; w_4_50<=Wgt_4_50; w_4_51<=Wgt_4_51; w_4_52<=Wgt_4_52; w_4_53<=Wgt_4_53; w_4_54<=Wgt_4_54; w_4_55<=Wgt_4_55; w_4_56<=Wgt_4_56; w_4_57<=Wgt_4_57; w_4_58<=Wgt_4_58; w_4_59<=Wgt_4_59; w_4_60<=Wgt_4_60; w_4_61<=Wgt_4_61; w_4_62<=Wgt_4_62; w_4_63<=Wgt_4_63; w_4_64<=Wgt_4_64; w_4_65<=Wgt_4_65; w_4_66<=Wgt_4_66; w_4_67<=Wgt_4_67; w_4_68<=Wgt_4_68; w_4_69<=Wgt_4_69; w_4_70<=Wgt_4_70; w_4_71<=Wgt_4_71; w_4_72<=Wgt_4_72; w_4_73<=Wgt_4_73; w_4_74<=Wgt_4_74; w_4_75<=Wgt_4_75; w_4_76<=Wgt_4_76; w_4_77<=Wgt_4_77; w_4_78<=Wgt_4_78; w_4_79<=Wgt_4_79; w_4_80<=Wgt_4_80; w_4_81<=Wgt_4_81; w_4_82<=Wgt_4_82; w_4_83<=Wgt_4_83; w_4_84<=Wgt_4_84; w_4_85<=Wgt_4_85; w_4_86<=Wgt_4_86; w_4_87<=Wgt_4_87; w_4_88<=Wgt_4_88; w_4_89<=Wgt_4_89; w_4_90<=Wgt_4_90; w_4_91<=Wgt_4_91; w_4_92<=Wgt_4_92; w_4_93<=Wgt_4_93; w_4_94<=Wgt_4_94; w_4_95<=Wgt_4_95; w_4_96<=Wgt_4_96; w_4_97<=Wgt_4_97; w_4_98<=Wgt_4_98; w_4_99<=Wgt_4_99; w_4_100<=Wgt_4_100; w_4_101<=Wgt_4_101; w_4_102<=Wgt_4_102; w_4_103<=Wgt_4_103; w_4_104<=Wgt_4_104; w_4_105<=Wgt_4_105; w_4_106<=Wgt_4_106; w_4_107<=Wgt_4_107; w_4_108<=Wgt_4_108; w_4_109<=Wgt_4_109; w_4_110<=Wgt_4_110; w_4_111<=Wgt_4_111; w_4_112<=Wgt_4_112; w_4_113<=Wgt_4_113; w_4_114<=Wgt_4_114; w_4_115<=Wgt_4_115; w_4_116<=Wgt_4_116; w_4_117<=Wgt_4_117; w_4_118<=Wgt_4_118; w_4_119<=Wgt_4_119; w_4_120<=Wgt_4_120; w_4_121<=Wgt_4_121; w_4_122<=Wgt_4_122; w_4_123<=Wgt_4_123; w_4_124<=Wgt_4_124; w_4_125<=Wgt_4_125; w_4_126<=Wgt_4_126; w_4_127<=Wgt_4_127; w_4_128<=Wgt_4_128; w_4_129<=Wgt_4_129; w_4_130<=Wgt_4_130; w_4_131<=Wgt_4_131; w_4_132<=Wgt_4_132; w_4_133<=Wgt_4_133; w_4_134<=Wgt_4_134; w_4_135<=Wgt_4_135; w_4_136<=Wgt_4_136; w_4_137<=Wgt_4_137; w_4_138<=Wgt_4_138; w_4_139<=Wgt_4_139; w_4_140<=Wgt_4_140; w_4_141<=Wgt_4_141; w_4_142<=Wgt_4_142; w_4_143<=Wgt_4_143; w_4_144<=Wgt_4_144; w_4_145<=Wgt_4_145; w_4_146<=Wgt_4_146; w_4_147<=Wgt_4_147; w_4_148<=Wgt_4_148; w_4_149<=Wgt_4_149; w_4_150<=Wgt_4_150; w_4_151<=Wgt_4_151; w_4_152<=Wgt_4_152; w_4_153<=Wgt_4_153; w_4_154<=Wgt_4_154; w_4_155<=Wgt_4_155; w_4_156<=Wgt_4_156; w_4_157<=Wgt_4_157; w_4_158<=Wgt_4_158; w_4_159<=Wgt_4_159; w_4_160<=Wgt_4_160; w_4_161<=Wgt_4_161; w_4_162<=Wgt_4_162; w_4_163<=Wgt_4_163; w_4_164<=Wgt_4_164; w_4_165<=Wgt_4_165; w_4_166<=Wgt_4_166; w_4_167<=Wgt_4_167; w_4_168<=Wgt_4_168; w_4_169<=Wgt_4_169; w_4_170<=Wgt_4_170; w_4_171<=Wgt_4_171; w_4_172<=Wgt_4_172; w_4_173<=Wgt_4_173; w_4_174<=Wgt_4_174; w_4_175<=Wgt_4_175; w_4_176<=Wgt_4_176; w_4_177<=Wgt_4_177; w_4_178<=Wgt_4_178; w_4_179<=Wgt_4_179; w_4_180<=Wgt_4_180; w_4_181<=Wgt_4_181; w_4_182<=Wgt_4_182; w_4_183<=Wgt_4_183; w_4_184<=Wgt_4_184; w_4_185<=Wgt_4_185; w_4_186<=Wgt_4_186; w_4_187<=Wgt_4_187; w_4_188<=Wgt_4_188; w_4_189<=Wgt_4_189; w_4_190<=Wgt_4_190; w_4_191<=Wgt_4_191; w_4_192<=Wgt_4_192; w_4_193<=Wgt_4_193; w_4_194<=Wgt_4_194; w_4_195<=Wgt_4_195; w_4_196<=Wgt_4_196; w_4_197<=Wgt_4_197; w_4_198<=Wgt_4_198; w_4_199<=Wgt_4_199; w_4_200<=Wgt_4_200; w_4_201<=Wgt_4_201; w_4_202<=Wgt_4_202; w_4_203<=Wgt_4_203; w_4_204<=Wgt_4_204; w_4_205<=Wgt_4_205; w_4_206<=Wgt_4_206; w_4_207<=Wgt_4_207; w_4_208<=Wgt_4_208; w_4_209<=Wgt_4_209; w_4_210<=Wgt_4_210; w_4_211<=Wgt_4_211; w_4_212<=Wgt_4_212; w_4_213<=Wgt_4_213; w_4_214<=Wgt_4_214; w_4_215<=Wgt_4_215; w_4_216<=Wgt_4_216; w_4_217<=Wgt_4_217; w_4_218<=Wgt_4_218; w_4_219<=Wgt_4_219; w_4_220<=Wgt_4_220; w_4_221<=Wgt_4_221; w_4_222<=Wgt_4_222; w_4_223<=Wgt_4_223; w_4_224<=Wgt_4_224; w_4_225<=Wgt_4_225; w_4_226<=Wgt_4_226; w_4_227<=Wgt_4_227; w_4_228<=Wgt_4_228; w_4_229<=Wgt_4_229; w_4_230<=Wgt_4_230; w_4_231<=Wgt_4_231; w_4_232<=Wgt_4_232; w_4_233<=Wgt_4_233; w_4_234<=Wgt_4_234; w_4_235<=Wgt_4_235; w_4_236<=Wgt_4_236; w_4_237<=Wgt_4_237; w_4_238<=Wgt_4_238; w_4_239<=Wgt_4_239; w_4_240<=Wgt_4_240; w_4_241<=Wgt_4_241; w_4_242<=Wgt_4_242; w_4_243<=Wgt_4_243; w_4_244<=Wgt_4_244; w_4_245<=Wgt_4_245; w_4_246<=Wgt_4_246; w_4_247<=Wgt_4_247; w_4_248<=Wgt_4_248; w_4_249<=Wgt_4_249; w_4_250<=Wgt_4_250; w_4_251<=Wgt_4_251; w_4_252<=Wgt_4_252; w_4_253<=Wgt_4_253; w_4_254<=Wgt_4_254; w_4_255<=Wgt_4_255; w_4_256<=Wgt_4_256; w_4_257<=Wgt_4_257; w_4_258<=Wgt_4_258; w_4_259<=Wgt_4_259; w_4_260<=Wgt_4_260; w_4_261<=Wgt_4_261; w_4_262<=Wgt_4_262; w_4_263<=Wgt_4_263; w_4_264<=Wgt_4_264; w_4_265<=Wgt_4_265; w_4_266<=Wgt_4_266; w_4_267<=Wgt_4_267; w_4_268<=Wgt_4_268; w_4_269<=Wgt_4_269; w_4_270<=Wgt_4_270; w_4_271<=Wgt_4_271; w_4_272<=Wgt_4_272; w_4_273<=Wgt_4_273; w_4_274<=Wgt_4_274; w_4_275<=Wgt_4_275; w_4_276<=Wgt_4_276; w_4_277<=Wgt_4_277; w_4_278<=Wgt_4_278; w_4_279<=Wgt_4_279; w_4_280<=Wgt_4_280; w_4_281<=Wgt_4_281; w_4_282<=Wgt_4_282; w_4_283<=Wgt_4_283; w_4_284<=Wgt_4_284; w_4_285<=Wgt_4_285; w_4_286<=Wgt_4_286; w_4_287<=Wgt_4_287; w_4_288<=Wgt_4_288; w_4_289<=Wgt_4_289; w_4_290<=Wgt_4_290; w_4_291<=Wgt_4_291; w_4_292<=Wgt_4_292; w_4_293<=Wgt_4_293; w_4_294<=Wgt_4_294; w_4_295<=Wgt_4_295; w_4_296<=Wgt_4_296; w_4_297<=Wgt_4_297; w_4_298<=Wgt_4_298; w_4_299<=Wgt_4_299; w_4_300<=Wgt_4_300; w_4_301<=Wgt_4_301; w_4_302<=Wgt_4_302; w_4_303<=Wgt_4_303; w_4_304<=Wgt_4_304; w_4_305<=Wgt_4_305; w_4_306<=Wgt_4_306; w_4_307<=Wgt_4_307; w_4_308<=Wgt_4_308; w_4_309<=Wgt_4_309; w_4_310<=Wgt_4_310; w_4_311<=Wgt_4_311; w_4_312<=Wgt_4_312; w_4_313<=Wgt_4_313; w_4_314<=Wgt_4_314; w_4_315<=Wgt_4_315; w_4_316<=Wgt_4_316; w_4_317<=Wgt_4_317; w_4_318<=Wgt_4_318; w_4_319<=Wgt_4_319; w_4_320<=Wgt_4_320; w_4_321<=Wgt_4_321; w_4_322<=Wgt_4_322; w_4_323<=Wgt_4_323; w_4_324<=Wgt_4_324; w_4_325<=Wgt_4_325; w_4_326<=Wgt_4_326; w_4_327<=Wgt_4_327; w_4_328<=Wgt_4_328; w_4_329<=Wgt_4_329; w_4_330<=Wgt_4_330; w_4_331<=Wgt_4_331; w_4_332<=Wgt_4_332; w_4_333<=Wgt_4_333; w_4_334<=Wgt_4_334; w_4_335<=Wgt_4_335; w_4_336<=Wgt_4_336; w_4_337<=Wgt_4_337; w_4_338<=Wgt_4_338; w_4_339<=Wgt_4_339; w_4_340<=Wgt_4_340; w_4_341<=Wgt_4_341; w_4_342<=Wgt_4_342; w_4_343<=Wgt_4_343; w_4_344<=Wgt_4_344; w_4_345<=Wgt_4_345; w_4_346<=Wgt_4_346; w_4_347<=Wgt_4_347; w_4_348<=Wgt_4_348; w_4_349<=Wgt_4_349; w_4_350<=Wgt_4_350; w_4_351<=Wgt_4_351; w_4_352<=Wgt_4_352; w_4_353<=Wgt_4_353; w_4_354<=Wgt_4_354; w_4_355<=Wgt_4_355; w_4_356<=Wgt_4_356; w_4_357<=Wgt_4_357; w_4_358<=Wgt_4_358; w_4_359<=Wgt_4_359; w_4_360<=Wgt_4_360; w_4_361<=Wgt_4_361; w_4_362<=Wgt_4_362; w_4_363<=Wgt_4_363; w_4_364<=Wgt_4_364; w_4_365<=Wgt_4_365; w_4_366<=Wgt_4_366; w_4_367<=Wgt_4_367; w_4_368<=Wgt_4_368; w_4_369<=Wgt_4_369; w_4_370<=Wgt_4_370; w_4_371<=Wgt_4_371; w_4_372<=Wgt_4_372; w_4_373<=Wgt_4_373; w_4_374<=Wgt_4_374; w_4_375<=Wgt_4_375; w_4_376<=Wgt_4_376; w_4_377<=Wgt_4_377; w_4_378<=Wgt_4_378; w_4_379<=Wgt_4_379; w_4_380<=Wgt_4_380; w_4_381<=Wgt_4_381; w_4_382<=Wgt_4_382; w_4_383<=Wgt_4_383; w_4_384<=Wgt_4_384; w_4_385<=Wgt_4_385; w_4_386<=Wgt_4_386; w_4_387<=Wgt_4_387; w_4_388<=Wgt_4_388; w_4_389<=Wgt_4_389; w_4_390<=Wgt_4_390; w_4_391<=Wgt_4_391; w_4_392<=Wgt_4_392; w_4_393<=Wgt_4_393; w_4_394<=Wgt_4_394; w_4_395<=Wgt_4_395; w_4_396<=Wgt_4_396; w_4_397<=Wgt_4_397; w_4_398<=Wgt_4_398; w_4_399<=Wgt_4_399; w_4_400<=Wgt_4_400; w_4_401<=Wgt_4_401; w_4_402<=Wgt_4_402; w_4_403<=Wgt_4_403; w_4_404<=Wgt_4_404; w_4_405<=Wgt_4_405; w_4_406<=Wgt_4_406; w_4_407<=Wgt_4_407; w_4_408<=Wgt_4_408; w_4_409<=Wgt_4_409; w_4_410<=Wgt_4_410; w_4_411<=Wgt_4_411; w_4_412<=Wgt_4_412; w_4_413<=Wgt_4_413; w_4_414<=Wgt_4_414; w_4_415<=Wgt_4_415; w_4_416<=Wgt_4_416; w_4_417<=Wgt_4_417; w_4_418<=Wgt_4_418; w_4_419<=Wgt_4_419; w_4_420<=Wgt_4_420; w_4_421<=Wgt_4_421; w_4_422<=Wgt_4_422; w_4_423<=Wgt_4_423; w_4_424<=Wgt_4_424; w_4_425<=Wgt_4_425; w_4_426<=Wgt_4_426; w_4_427<=Wgt_4_427; w_4_428<=Wgt_4_428; w_4_429<=Wgt_4_429; w_4_430<=Wgt_4_430; w_4_431<=Wgt_4_431; w_4_432<=Wgt_4_432; w_4_433<=Wgt_4_433; w_4_434<=Wgt_4_434; w_4_435<=Wgt_4_435; w_4_436<=Wgt_4_436; w_4_437<=Wgt_4_437; w_4_438<=Wgt_4_438; w_4_439<=Wgt_4_439; w_4_440<=Wgt_4_440; w_4_441<=Wgt_4_441; w_4_442<=Wgt_4_442; w_4_443<=Wgt_4_443; w_4_444<=Wgt_4_444; w_4_445<=Wgt_4_445; w_4_446<=Wgt_4_446; w_4_447<=Wgt_4_447; w_4_448<=Wgt_4_448; w_4_449<=Wgt_4_449; w_4_450<=Wgt_4_450; w_4_451<=Wgt_4_451; w_4_452<=Wgt_4_452; w_4_453<=Wgt_4_453; w_4_454<=Wgt_4_454; w_4_455<=Wgt_4_455; w_4_456<=Wgt_4_456; w_4_457<=Wgt_4_457; w_4_458<=Wgt_4_458; w_4_459<=Wgt_4_459; w_4_460<=Wgt_4_460; w_4_461<=Wgt_4_461; w_4_462<=Wgt_4_462; w_4_463<=Wgt_4_463; w_4_464<=Wgt_4_464; w_4_465<=Wgt_4_465; w_4_466<=Wgt_4_466; w_4_467<=Wgt_4_467; w_4_468<=Wgt_4_468; w_4_469<=Wgt_4_469; w_4_470<=Wgt_4_470; w_4_471<=Wgt_4_471; w_4_472<=Wgt_4_472; w_4_473<=Wgt_4_473; w_4_474<=Wgt_4_474; w_4_475<=Wgt_4_475; w_4_476<=Wgt_4_476; w_4_477<=Wgt_4_477; w_4_478<=Wgt_4_478; w_4_479<=Wgt_4_479; w_4_480<=Wgt_4_480; w_4_481<=Wgt_4_481; w_4_482<=Wgt_4_482; w_4_483<=Wgt_4_483; w_4_484<=Wgt_4_484; w_4_485<=Wgt_4_485; w_4_486<=Wgt_4_486; w_4_487<=Wgt_4_487; w_4_488<=Wgt_4_488; w_4_489<=Wgt_4_489; w_4_490<=Wgt_4_490; w_4_491<=Wgt_4_491; w_4_492<=Wgt_4_492; w_4_493<=Wgt_4_493; w_4_494<=Wgt_4_494; w_4_495<=Wgt_4_495; w_4_496<=Wgt_4_496; w_4_497<=Wgt_4_497; w_4_498<=Wgt_4_498; w_4_499<=Wgt_4_499; w_4_500<=Wgt_4_500; w_4_501<=Wgt_4_501; w_4_502<=Wgt_4_502; w_4_503<=Wgt_4_503; w_4_504<=Wgt_4_504; w_4_505<=Wgt_4_505; w_4_506<=Wgt_4_506; w_4_507<=Wgt_4_507; w_4_508<=Wgt_4_508; w_4_509<=Wgt_4_509; w_4_510<=Wgt_4_510; w_4_511<=Wgt_4_511; w_4_512<=Wgt_4_512; w_4_513<=Wgt_4_513; w_4_514<=Wgt_4_514; w_4_515<=Wgt_4_515; w_4_516<=Wgt_4_516; w_4_517<=Wgt_4_517; w_4_518<=Wgt_4_518; w_4_519<=Wgt_4_519; w_4_520<=Wgt_4_520; w_4_521<=Wgt_4_521; w_4_522<=Wgt_4_522; w_4_523<=Wgt_4_523; w_4_524<=Wgt_4_524; w_4_525<=Wgt_4_525; w_4_526<=Wgt_4_526; w_4_527<=Wgt_4_527; w_4_528<=Wgt_4_528; w_4_529<=Wgt_4_529; w_4_530<=Wgt_4_530; w_4_531<=Wgt_4_531; w_4_532<=Wgt_4_532; w_4_533<=Wgt_4_533; w_4_534<=Wgt_4_534; w_4_535<=Wgt_4_535; w_4_536<=Wgt_4_536; w_4_537<=Wgt_4_537; w_4_538<=Wgt_4_538; w_4_539<=Wgt_4_539; w_4_540<=Wgt_4_540; w_4_541<=Wgt_4_541; w_4_542<=Wgt_4_542; w_4_543<=Wgt_4_543; w_4_544<=Wgt_4_544; w_4_545<=Wgt_4_545; w_4_546<=Wgt_4_546; w_4_547<=Wgt_4_547; w_4_548<=Wgt_4_548; w_4_549<=Wgt_4_549; w_4_550<=Wgt_4_550; w_4_551<=Wgt_4_551; w_4_552<=Wgt_4_552; w_4_553<=Wgt_4_553; w_4_554<=Wgt_4_554; w_4_555<=Wgt_4_555; w_4_556<=Wgt_4_556; w_4_557<=Wgt_4_557; w_4_558<=Wgt_4_558; w_4_559<=Wgt_4_559; w_4_560<=Wgt_4_560; w_4_561<=Wgt_4_561; w_4_562<=Wgt_4_562; w_4_563<=Wgt_4_563; w_4_564<=Wgt_4_564; w_4_565<=Wgt_4_565; w_4_566<=Wgt_4_566; w_4_567<=Wgt_4_567; w_4_568<=Wgt_4_568; w_4_569<=Wgt_4_569; w_4_570<=Wgt_4_570; w_4_571<=Wgt_4_571; w_4_572<=Wgt_4_572; w_4_573<=Wgt_4_573; w_4_574<=Wgt_4_574; w_4_575<=Wgt_4_575; w_4_576<=Wgt_4_576; w_4_577<=Wgt_4_577; w_4_578<=Wgt_4_578; w_4_579<=Wgt_4_579; w_4_580<=Wgt_4_580; w_4_581<=Wgt_4_581; w_4_582<=Wgt_4_582; w_4_583<=Wgt_4_583; w_4_584<=Wgt_4_584; w_4_585<=Wgt_4_585; w_4_586<=Wgt_4_586; w_4_587<=Wgt_4_587; w_4_588<=Wgt_4_588; w_4_589<=Wgt_4_589; w_4_590<=Wgt_4_590; w_4_591<=Wgt_4_591; w_4_592<=Wgt_4_592; w_4_593<=Wgt_4_593; w_4_594<=Wgt_4_594; w_4_595<=Wgt_4_595; w_4_596<=Wgt_4_596; w_4_597<=Wgt_4_597; w_4_598<=Wgt_4_598; w_4_599<=Wgt_4_599; w_4_600<=Wgt_4_600; w_4_601<=Wgt_4_601; w_4_602<=Wgt_4_602; w_4_603<=Wgt_4_603; w_4_604<=Wgt_4_604; w_4_605<=Wgt_4_605; w_4_606<=Wgt_4_606; w_4_607<=Wgt_4_607; w_4_608<=Wgt_4_608; w_4_609<=Wgt_4_609; w_4_610<=Wgt_4_610; w_4_611<=Wgt_4_611; w_4_612<=Wgt_4_612; w_4_613<=Wgt_4_613; w_4_614<=Wgt_4_614; w_4_615<=Wgt_4_615; w_4_616<=Wgt_4_616; w_4_617<=Wgt_4_617; w_4_618<=Wgt_4_618; w_4_619<=Wgt_4_619; w_4_620<=Wgt_4_620; w_4_621<=Wgt_4_621; w_4_622<=Wgt_4_622; w_4_623<=Wgt_4_623; w_4_624<=Wgt_4_624; w_4_625<=Wgt_4_625; w_4_626<=Wgt_4_626; w_4_627<=Wgt_4_627; w_4_628<=Wgt_4_628; w_4_629<=Wgt_4_629; w_4_630<=Wgt_4_630; w_4_631<=Wgt_4_631; w_4_632<=Wgt_4_632; w_4_633<=Wgt_4_633; w_4_634<=Wgt_4_634; w_4_635<=Wgt_4_635; w_4_636<=Wgt_4_636; w_4_637<=Wgt_4_637; w_4_638<=Wgt_4_638; w_4_639<=Wgt_4_639; w_4_640<=Wgt_4_640; w_4_641<=Wgt_4_641; w_4_642<=Wgt_4_642; w_4_643<=Wgt_4_643; w_4_644<=Wgt_4_644; w_4_645<=Wgt_4_645; w_4_646<=Wgt_4_646; w_4_647<=Wgt_4_647; w_4_648<=Wgt_4_648; w_4_649<=Wgt_4_649; w_4_650<=Wgt_4_650; w_4_651<=Wgt_4_651; w_4_652<=Wgt_4_652; w_4_653<=Wgt_4_653; w_4_654<=Wgt_4_654; w_4_655<=Wgt_4_655; w_4_656<=Wgt_4_656; w_4_657<=Wgt_4_657; w_4_658<=Wgt_4_658; w_4_659<=Wgt_4_659; w_4_660<=Wgt_4_660; w_4_661<=Wgt_4_661; w_4_662<=Wgt_4_662; w_4_663<=Wgt_4_663; w_4_664<=Wgt_4_664; w_4_665<=Wgt_4_665; w_4_666<=Wgt_4_666; w_4_667<=Wgt_4_667; w_4_668<=Wgt_4_668; w_4_669<=Wgt_4_669; w_4_670<=Wgt_4_670; w_4_671<=Wgt_4_671; w_4_672<=Wgt_4_672; w_4_673<=Wgt_4_673; w_4_674<=Wgt_4_674; w_4_675<=Wgt_4_675; w_4_676<=Wgt_4_676; w_4_677<=Wgt_4_677; w_4_678<=Wgt_4_678; w_4_679<=Wgt_4_679; w_4_680<=Wgt_4_680; w_4_681<=Wgt_4_681; w_4_682<=Wgt_4_682; w_4_683<=Wgt_4_683; w_4_684<=Wgt_4_684; w_4_685<=Wgt_4_685; w_4_686<=Wgt_4_686; w_4_687<=Wgt_4_687; w_4_688<=Wgt_4_688; w_4_689<=Wgt_4_689; w_4_690<=Wgt_4_690; w_4_691<=Wgt_4_691; w_4_692<=Wgt_4_692; w_4_693<=Wgt_4_693; w_4_694<=Wgt_4_694; w_4_695<=Wgt_4_695; w_4_696<=Wgt_4_696; w_4_697<=Wgt_4_697; w_4_698<=Wgt_4_698; w_4_699<=Wgt_4_699; w_4_700<=Wgt_4_700; w_4_701<=Wgt_4_701; w_4_702<=Wgt_4_702; w_4_703<=Wgt_4_703; w_4_704<=Wgt_4_704; w_4_705<=Wgt_4_705; w_4_706<=Wgt_4_706; w_4_707<=Wgt_4_707; w_4_708<=Wgt_4_708; w_4_709<=Wgt_4_709; w_4_710<=Wgt_4_710; w_4_711<=Wgt_4_711; w_4_712<=Wgt_4_712; w_4_713<=Wgt_4_713; w_4_714<=Wgt_4_714; w_4_715<=Wgt_4_715; w_4_716<=Wgt_4_716; w_4_717<=Wgt_4_717; w_4_718<=Wgt_4_718; w_4_719<=Wgt_4_719; w_4_720<=Wgt_4_720; w_4_721<=Wgt_4_721; w_4_722<=Wgt_4_722; w_4_723<=Wgt_4_723; w_4_724<=Wgt_4_724; w_4_725<=Wgt_4_725; w_4_726<=Wgt_4_726; w_4_727<=Wgt_4_727; w_4_728<=Wgt_4_728; w_4_729<=Wgt_4_729; w_4_730<=Wgt_4_730; w_4_731<=Wgt_4_731; w_4_732<=Wgt_4_732; w_4_733<=Wgt_4_733; w_4_734<=Wgt_4_734; w_4_735<=Wgt_4_735; w_4_736<=Wgt_4_736; w_4_737<=Wgt_4_737; w_4_738<=Wgt_4_738; w_4_739<=Wgt_4_739; w_4_740<=Wgt_4_740; w_4_741<=Wgt_4_741; w_4_742<=Wgt_4_742; w_4_743<=Wgt_4_743; w_4_744<=Wgt_4_744; w_4_745<=Wgt_4_745; w_4_746<=Wgt_4_746; w_4_747<=Wgt_4_747; w_4_748<=Wgt_4_748; w_4_749<=Wgt_4_749; w_4_750<=Wgt_4_750; w_4_751<=Wgt_4_751; w_4_752<=Wgt_4_752; w_4_753<=Wgt_4_753; w_4_754<=Wgt_4_754; w_4_755<=Wgt_4_755; w_4_756<=Wgt_4_756; w_4_757<=Wgt_4_757; w_4_758<=Wgt_4_758; w_4_759<=Wgt_4_759; w_4_760<=Wgt_4_760; w_4_761<=Wgt_4_761; w_4_762<=Wgt_4_762; w_4_763<=Wgt_4_763; w_4_764<=Wgt_4_764; w_4_765<=Wgt_4_765; w_4_766<=Wgt_4_766; w_4_767<=Wgt_4_767; w_4_768<=Wgt_4_768; w_4_769<=Wgt_4_769; w_4_770<=Wgt_4_770; w_4_771<=Wgt_4_771; w_4_772<=Wgt_4_772; w_4_773<=Wgt_4_773; w_4_774<=Wgt_4_774; w_4_775<=Wgt_4_775; w_4_776<=Wgt_4_776; w_4_777<=Wgt_4_777; w_4_778<=Wgt_4_778; w_4_779<=Wgt_4_779; w_4_780<=Wgt_4_780; w_4_781<=Wgt_4_781; w_4_782<=Wgt_4_782; w_4_783<=Wgt_4_783; w_4_784<=Wgt_4_784; 
					w_5_0<=Wgt_5_0; w_5_1<=Wgt_5_1; w_5_2<=Wgt_5_2; w_5_3<=Wgt_5_3; w_5_4<=Wgt_5_4; w_5_5<=Wgt_5_5; w_5_6<=Wgt_5_6; w_5_7<=Wgt_5_7; w_5_8<=Wgt_5_8; w_5_9<=Wgt_5_9; w_5_10<=Wgt_5_10; w_5_11<=Wgt_5_11; w_5_12<=Wgt_5_12; w_5_13<=Wgt_5_13; w_5_14<=Wgt_5_14; w_5_15<=Wgt_5_15; w_5_16<=Wgt_5_16; w_5_17<=Wgt_5_17; w_5_18<=Wgt_5_18; w_5_19<=Wgt_5_19; w_5_20<=Wgt_5_20; w_5_21<=Wgt_5_21; w_5_22<=Wgt_5_22; w_5_23<=Wgt_5_23; w_5_24<=Wgt_5_24; w_5_25<=Wgt_5_25; w_5_26<=Wgt_5_26; w_5_27<=Wgt_5_27; w_5_28<=Wgt_5_28; w_5_29<=Wgt_5_29; w_5_30<=Wgt_5_30; w_5_31<=Wgt_5_31; w_5_32<=Wgt_5_32; w_5_33<=Wgt_5_33; w_5_34<=Wgt_5_34; w_5_35<=Wgt_5_35; w_5_36<=Wgt_5_36; w_5_37<=Wgt_5_37; w_5_38<=Wgt_5_38; w_5_39<=Wgt_5_39; w_5_40<=Wgt_5_40; w_5_41<=Wgt_5_41; w_5_42<=Wgt_5_42; w_5_43<=Wgt_5_43; w_5_44<=Wgt_5_44; w_5_45<=Wgt_5_45; w_5_46<=Wgt_5_46; w_5_47<=Wgt_5_47; w_5_48<=Wgt_5_48; w_5_49<=Wgt_5_49; w_5_50<=Wgt_5_50; w_5_51<=Wgt_5_51; w_5_52<=Wgt_5_52; w_5_53<=Wgt_5_53; w_5_54<=Wgt_5_54; w_5_55<=Wgt_5_55; w_5_56<=Wgt_5_56; w_5_57<=Wgt_5_57; w_5_58<=Wgt_5_58; w_5_59<=Wgt_5_59; w_5_60<=Wgt_5_60; w_5_61<=Wgt_5_61; w_5_62<=Wgt_5_62; w_5_63<=Wgt_5_63; w_5_64<=Wgt_5_64; w_5_65<=Wgt_5_65; w_5_66<=Wgt_5_66; w_5_67<=Wgt_5_67; w_5_68<=Wgt_5_68; w_5_69<=Wgt_5_69; w_5_70<=Wgt_5_70; w_5_71<=Wgt_5_71; w_5_72<=Wgt_5_72; w_5_73<=Wgt_5_73; w_5_74<=Wgt_5_74; w_5_75<=Wgt_5_75; w_5_76<=Wgt_5_76; w_5_77<=Wgt_5_77; w_5_78<=Wgt_5_78; w_5_79<=Wgt_5_79; w_5_80<=Wgt_5_80; w_5_81<=Wgt_5_81; w_5_82<=Wgt_5_82; w_5_83<=Wgt_5_83; w_5_84<=Wgt_5_84; w_5_85<=Wgt_5_85; w_5_86<=Wgt_5_86; w_5_87<=Wgt_5_87; w_5_88<=Wgt_5_88; w_5_89<=Wgt_5_89; w_5_90<=Wgt_5_90; w_5_91<=Wgt_5_91; w_5_92<=Wgt_5_92; w_5_93<=Wgt_5_93; w_5_94<=Wgt_5_94; w_5_95<=Wgt_5_95; w_5_96<=Wgt_5_96; w_5_97<=Wgt_5_97; w_5_98<=Wgt_5_98; w_5_99<=Wgt_5_99; w_5_100<=Wgt_5_100; w_5_101<=Wgt_5_101; w_5_102<=Wgt_5_102; w_5_103<=Wgt_5_103; w_5_104<=Wgt_5_104; w_5_105<=Wgt_5_105; w_5_106<=Wgt_5_106; w_5_107<=Wgt_5_107; w_5_108<=Wgt_5_108; w_5_109<=Wgt_5_109; w_5_110<=Wgt_5_110; w_5_111<=Wgt_5_111; w_5_112<=Wgt_5_112; w_5_113<=Wgt_5_113; w_5_114<=Wgt_5_114; w_5_115<=Wgt_5_115; w_5_116<=Wgt_5_116; w_5_117<=Wgt_5_117; w_5_118<=Wgt_5_118; w_5_119<=Wgt_5_119; w_5_120<=Wgt_5_120; w_5_121<=Wgt_5_121; w_5_122<=Wgt_5_122; w_5_123<=Wgt_5_123; w_5_124<=Wgt_5_124; w_5_125<=Wgt_5_125; w_5_126<=Wgt_5_126; w_5_127<=Wgt_5_127; w_5_128<=Wgt_5_128; w_5_129<=Wgt_5_129; w_5_130<=Wgt_5_130; w_5_131<=Wgt_5_131; w_5_132<=Wgt_5_132; w_5_133<=Wgt_5_133; w_5_134<=Wgt_5_134; w_5_135<=Wgt_5_135; w_5_136<=Wgt_5_136; w_5_137<=Wgt_5_137; w_5_138<=Wgt_5_138; w_5_139<=Wgt_5_139; w_5_140<=Wgt_5_140; w_5_141<=Wgt_5_141; w_5_142<=Wgt_5_142; w_5_143<=Wgt_5_143; w_5_144<=Wgt_5_144; w_5_145<=Wgt_5_145; w_5_146<=Wgt_5_146; w_5_147<=Wgt_5_147; w_5_148<=Wgt_5_148; w_5_149<=Wgt_5_149; w_5_150<=Wgt_5_150; w_5_151<=Wgt_5_151; w_5_152<=Wgt_5_152; w_5_153<=Wgt_5_153; w_5_154<=Wgt_5_154; w_5_155<=Wgt_5_155; w_5_156<=Wgt_5_156; w_5_157<=Wgt_5_157; w_5_158<=Wgt_5_158; w_5_159<=Wgt_5_159; w_5_160<=Wgt_5_160; w_5_161<=Wgt_5_161; w_5_162<=Wgt_5_162; w_5_163<=Wgt_5_163; w_5_164<=Wgt_5_164; w_5_165<=Wgt_5_165; w_5_166<=Wgt_5_166; w_5_167<=Wgt_5_167; w_5_168<=Wgt_5_168; w_5_169<=Wgt_5_169; w_5_170<=Wgt_5_170; w_5_171<=Wgt_5_171; w_5_172<=Wgt_5_172; w_5_173<=Wgt_5_173; w_5_174<=Wgt_5_174; w_5_175<=Wgt_5_175; w_5_176<=Wgt_5_176; w_5_177<=Wgt_5_177; w_5_178<=Wgt_5_178; w_5_179<=Wgt_5_179; w_5_180<=Wgt_5_180; w_5_181<=Wgt_5_181; w_5_182<=Wgt_5_182; w_5_183<=Wgt_5_183; w_5_184<=Wgt_5_184; w_5_185<=Wgt_5_185; w_5_186<=Wgt_5_186; w_5_187<=Wgt_5_187; w_5_188<=Wgt_5_188; w_5_189<=Wgt_5_189; w_5_190<=Wgt_5_190; w_5_191<=Wgt_5_191; w_5_192<=Wgt_5_192; w_5_193<=Wgt_5_193; w_5_194<=Wgt_5_194; w_5_195<=Wgt_5_195; w_5_196<=Wgt_5_196; w_5_197<=Wgt_5_197; w_5_198<=Wgt_5_198; w_5_199<=Wgt_5_199; w_5_200<=Wgt_5_200; w_5_201<=Wgt_5_201; w_5_202<=Wgt_5_202; w_5_203<=Wgt_5_203; w_5_204<=Wgt_5_204; w_5_205<=Wgt_5_205; w_5_206<=Wgt_5_206; w_5_207<=Wgt_5_207; w_5_208<=Wgt_5_208; w_5_209<=Wgt_5_209; w_5_210<=Wgt_5_210; w_5_211<=Wgt_5_211; w_5_212<=Wgt_5_212; w_5_213<=Wgt_5_213; w_5_214<=Wgt_5_214; w_5_215<=Wgt_5_215; w_5_216<=Wgt_5_216; w_5_217<=Wgt_5_217; w_5_218<=Wgt_5_218; w_5_219<=Wgt_5_219; w_5_220<=Wgt_5_220; w_5_221<=Wgt_5_221; w_5_222<=Wgt_5_222; w_5_223<=Wgt_5_223; w_5_224<=Wgt_5_224; w_5_225<=Wgt_5_225; w_5_226<=Wgt_5_226; w_5_227<=Wgt_5_227; w_5_228<=Wgt_5_228; w_5_229<=Wgt_5_229; w_5_230<=Wgt_5_230; w_5_231<=Wgt_5_231; w_5_232<=Wgt_5_232; w_5_233<=Wgt_5_233; w_5_234<=Wgt_5_234; w_5_235<=Wgt_5_235; w_5_236<=Wgt_5_236; w_5_237<=Wgt_5_237; w_5_238<=Wgt_5_238; w_5_239<=Wgt_5_239; w_5_240<=Wgt_5_240; w_5_241<=Wgt_5_241; w_5_242<=Wgt_5_242; w_5_243<=Wgt_5_243; w_5_244<=Wgt_5_244; w_5_245<=Wgt_5_245; w_5_246<=Wgt_5_246; w_5_247<=Wgt_5_247; w_5_248<=Wgt_5_248; w_5_249<=Wgt_5_249; w_5_250<=Wgt_5_250; w_5_251<=Wgt_5_251; w_5_252<=Wgt_5_252; w_5_253<=Wgt_5_253; w_5_254<=Wgt_5_254; w_5_255<=Wgt_5_255; w_5_256<=Wgt_5_256; w_5_257<=Wgt_5_257; w_5_258<=Wgt_5_258; w_5_259<=Wgt_5_259; w_5_260<=Wgt_5_260; w_5_261<=Wgt_5_261; w_5_262<=Wgt_5_262; w_5_263<=Wgt_5_263; w_5_264<=Wgt_5_264; w_5_265<=Wgt_5_265; w_5_266<=Wgt_5_266; w_5_267<=Wgt_5_267; w_5_268<=Wgt_5_268; w_5_269<=Wgt_5_269; w_5_270<=Wgt_5_270; w_5_271<=Wgt_5_271; w_5_272<=Wgt_5_272; w_5_273<=Wgt_5_273; w_5_274<=Wgt_5_274; w_5_275<=Wgt_5_275; w_5_276<=Wgt_5_276; w_5_277<=Wgt_5_277; w_5_278<=Wgt_5_278; w_5_279<=Wgt_5_279; w_5_280<=Wgt_5_280; w_5_281<=Wgt_5_281; w_5_282<=Wgt_5_282; w_5_283<=Wgt_5_283; w_5_284<=Wgt_5_284; w_5_285<=Wgt_5_285; w_5_286<=Wgt_5_286; w_5_287<=Wgt_5_287; w_5_288<=Wgt_5_288; w_5_289<=Wgt_5_289; w_5_290<=Wgt_5_290; w_5_291<=Wgt_5_291; w_5_292<=Wgt_5_292; w_5_293<=Wgt_5_293; w_5_294<=Wgt_5_294; w_5_295<=Wgt_5_295; w_5_296<=Wgt_5_296; w_5_297<=Wgt_5_297; w_5_298<=Wgt_5_298; w_5_299<=Wgt_5_299; w_5_300<=Wgt_5_300; w_5_301<=Wgt_5_301; w_5_302<=Wgt_5_302; w_5_303<=Wgt_5_303; w_5_304<=Wgt_5_304; w_5_305<=Wgt_5_305; w_5_306<=Wgt_5_306; w_5_307<=Wgt_5_307; w_5_308<=Wgt_5_308; w_5_309<=Wgt_5_309; w_5_310<=Wgt_5_310; w_5_311<=Wgt_5_311; w_5_312<=Wgt_5_312; w_5_313<=Wgt_5_313; w_5_314<=Wgt_5_314; w_5_315<=Wgt_5_315; w_5_316<=Wgt_5_316; w_5_317<=Wgt_5_317; w_5_318<=Wgt_5_318; w_5_319<=Wgt_5_319; w_5_320<=Wgt_5_320; w_5_321<=Wgt_5_321; w_5_322<=Wgt_5_322; w_5_323<=Wgt_5_323; w_5_324<=Wgt_5_324; w_5_325<=Wgt_5_325; w_5_326<=Wgt_5_326; w_5_327<=Wgt_5_327; w_5_328<=Wgt_5_328; w_5_329<=Wgt_5_329; w_5_330<=Wgt_5_330; w_5_331<=Wgt_5_331; w_5_332<=Wgt_5_332; w_5_333<=Wgt_5_333; w_5_334<=Wgt_5_334; w_5_335<=Wgt_5_335; w_5_336<=Wgt_5_336; w_5_337<=Wgt_5_337; w_5_338<=Wgt_5_338; w_5_339<=Wgt_5_339; w_5_340<=Wgt_5_340; w_5_341<=Wgt_5_341; w_5_342<=Wgt_5_342; w_5_343<=Wgt_5_343; w_5_344<=Wgt_5_344; w_5_345<=Wgt_5_345; w_5_346<=Wgt_5_346; w_5_347<=Wgt_5_347; w_5_348<=Wgt_5_348; w_5_349<=Wgt_5_349; w_5_350<=Wgt_5_350; w_5_351<=Wgt_5_351; w_5_352<=Wgt_5_352; w_5_353<=Wgt_5_353; w_5_354<=Wgt_5_354; w_5_355<=Wgt_5_355; w_5_356<=Wgt_5_356; w_5_357<=Wgt_5_357; w_5_358<=Wgt_5_358; w_5_359<=Wgt_5_359; w_5_360<=Wgt_5_360; w_5_361<=Wgt_5_361; w_5_362<=Wgt_5_362; w_5_363<=Wgt_5_363; w_5_364<=Wgt_5_364; w_5_365<=Wgt_5_365; w_5_366<=Wgt_5_366; w_5_367<=Wgt_5_367; w_5_368<=Wgt_5_368; w_5_369<=Wgt_5_369; w_5_370<=Wgt_5_370; w_5_371<=Wgt_5_371; w_5_372<=Wgt_5_372; w_5_373<=Wgt_5_373; w_5_374<=Wgt_5_374; w_5_375<=Wgt_5_375; w_5_376<=Wgt_5_376; w_5_377<=Wgt_5_377; w_5_378<=Wgt_5_378; w_5_379<=Wgt_5_379; w_5_380<=Wgt_5_380; w_5_381<=Wgt_5_381; w_5_382<=Wgt_5_382; w_5_383<=Wgt_5_383; w_5_384<=Wgt_5_384; w_5_385<=Wgt_5_385; w_5_386<=Wgt_5_386; w_5_387<=Wgt_5_387; w_5_388<=Wgt_5_388; w_5_389<=Wgt_5_389; w_5_390<=Wgt_5_390; w_5_391<=Wgt_5_391; w_5_392<=Wgt_5_392; w_5_393<=Wgt_5_393; w_5_394<=Wgt_5_394; w_5_395<=Wgt_5_395; w_5_396<=Wgt_5_396; w_5_397<=Wgt_5_397; w_5_398<=Wgt_5_398; w_5_399<=Wgt_5_399; w_5_400<=Wgt_5_400; w_5_401<=Wgt_5_401; w_5_402<=Wgt_5_402; w_5_403<=Wgt_5_403; w_5_404<=Wgt_5_404; w_5_405<=Wgt_5_405; w_5_406<=Wgt_5_406; w_5_407<=Wgt_5_407; w_5_408<=Wgt_5_408; w_5_409<=Wgt_5_409; w_5_410<=Wgt_5_410; w_5_411<=Wgt_5_411; w_5_412<=Wgt_5_412; w_5_413<=Wgt_5_413; w_5_414<=Wgt_5_414; w_5_415<=Wgt_5_415; w_5_416<=Wgt_5_416; w_5_417<=Wgt_5_417; w_5_418<=Wgt_5_418; w_5_419<=Wgt_5_419; w_5_420<=Wgt_5_420; w_5_421<=Wgt_5_421; w_5_422<=Wgt_5_422; w_5_423<=Wgt_5_423; w_5_424<=Wgt_5_424; w_5_425<=Wgt_5_425; w_5_426<=Wgt_5_426; w_5_427<=Wgt_5_427; w_5_428<=Wgt_5_428; w_5_429<=Wgt_5_429; w_5_430<=Wgt_5_430; w_5_431<=Wgt_5_431; w_5_432<=Wgt_5_432; w_5_433<=Wgt_5_433; w_5_434<=Wgt_5_434; w_5_435<=Wgt_5_435; w_5_436<=Wgt_5_436; w_5_437<=Wgt_5_437; w_5_438<=Wgt_5_438; w_5_439<=Wgt_5_439; w_5_440<=Wgt_5_440; w_5_441<=Wgt_5_441; w_5_442<=Wgt_5_442; w_5_443<=Wgt_5_443; w_5_444<=Wgt_5_444; w_5_445<=Wgt_5_445; w_5_446<=Wgt_5_446; w_5_447<=Wgt_5_447; w_5_448<=Wgt_5_448; w_5_449<=Wgt_5_449; w_5_450<=Wgt_5_450; w_5_451<=Wgt_5_451; w_5_452<=Wgt_5_452; w_5_453<=Wgt_5_453; w_5_454<=Wgt_5_454; w_5_455<=Wgt_5_455; w_5_456<=Wgt_5_456; w_5_457<=Wgt_5_457; w_5_458<=Wgt_5_458; w_5_459<=Wgt_5_459; w_5_460<=Wgt_5_460; w_5_461<=Wgt_5_461; w_5_462<=Wgt_5_462; w_5_463<=Wgt_5_463; w_5_464<=Wgt_5_464; w_5_465<=Wgt_5_465; w_5_466<=Wgt_5_466; w_5_467<=Wgt_5_467; w_5_468<=Wgt_5_468; w_5_469<=Wgt_5_469; w_5_470<=Wgt_5_470; w_5_471<=Wgt_5_471; w_5_472<=Wgt_5_472; w_5_473<=Wgt_5_473; w_5_474<=Wgt_5_474; w_5_475<=Wgt_5_475; w_5_476<=Wgt_5_476; w_5_477<=Wgt_5_477; w_5_478<=Wgt_5_478; w_5_479<=Wgt_5_479; w_5_480<=Wgt_5_480; w_5_481<=Wgt_5_481; w_5_482<=Wgt_5_482; w_5_483<=Wgt_5_483; w_5_484<=Wgt_5_484; w_5_485<=Wgt_5_485; w_5_486<=Wgt_5_486; w_5_487<=Wgt_5_487; w_5_488<=Wgt_5_488; w_5_489<=Wgt_5_489; w_5_490<=Wgt_5_490; w_5_491<=Wgt_5_491; w_5_492<=Wgt_5_492; w_5_493<=Wgt_5_493; w_5_494<=Wgt_5_494; w_5_495<=Wgt_5_495; w_5_496<=Wgt_5_496; w_5_497<=Wgt_5_497; w_5_498<=Wgt_5_498; w_5_499<=Wgt_5_499; w_5_500<=Wgt_5_500; w_5_501<=Wgt_5_501; w_5_502<=Wgt_5_502; w_5_503<=Wgt_5_503; w_5_504<=Wgt_5_504; w_5_505<=Wgt_5_505; w_5_506<=Wgt_5_506; w_5_507<=Wgt_5_507; w_5_508<=Wgt_5_508; w_5_509<=Wgt_5_509; w_5_510<=Wgt_5_510; w_5_511<=Wgt_5_511; w_5_512<=Wgt_5_512; w_5_513<=Wgt_5_513; w_5_514<=Wgt_5_514; w_5_515<=Wgt_5_515; w_5_516<=Wgt_5_516; w_5_517<=Wgt_5_517; w_5_518<=Wgt_5_518; w_5_519<=Wgt_5_519; w_5_520<=Wgt_5_520; w_5_521<=Wgt_5_521; w_5_522<=Wgt_5_522; w_5_523<=Wgt_5_523; w_5_524<=Wgt_5_524; w_5_525<=Wgt_5_525; w_5_526<=Wgt_5_526; w_5_527<=Wgt_5_527; w_5_528<=Wgt_5_528; w_5_529<=Wgt_5_529; w_5_530<=Wgt_5_530; w_5_531<=Wgt_5_531; w_5_532<=Wgt_5_532; w_5_533<=Wgt_5_533; w_5_534<=Wgt_5_534; w_5_535<=Wgt_5_535; w_5_536<=Wgt_5_536; w_5_537<=Wgt_5_537; w_5_538<=Wgt_5_538; w_5_539<=Wgt_5_539; w_5_540<=Wgt_5_540; w_5_541<=Wgt_5_541; w_5_542<=Wgt_5_542; w_5_543<=Wgt_5_543; w_5_544<=Wgt_5_544; w_5_545<=Wgt_5_545; w_5_546<=Wgt_5_546; w_5_547<=Wgt_5_547; w_5_548<=Wgt_5_548; w_5_549<=Wgt_5_549; w_5_550<=Wgt_5_550; w_5_551<=Wgt_5_551; w_5_552<=Wgt_5_552; w_5_553<=Wgt_5_553; w_5_554<=Wgt_5_554; w_5_555<=Wgt_5_555; w_5_556<=Wgt_5_556; w_5_557<=Wgt_5_557; w_5_558<=Wgt_5_558; w_5_559<=Wgt_5_559; w_5_560<=Wgt_5_560; w_5_561<=Wgt_5_561; w_5_562<=Wgt_5_562; w_5_563<=Wgt_5_563; w_5_564<=Wgt_5_564; w_5_565<=Wgt_5_565; w_5_566<=Wgt_5_566; w_5_567<=Wgt_5_567; w_5_568<=Wgt_5_568; w_5_569<=Wgt_5_569; w_5_570<=Wgt_5_570; w_5_571<=Wgt_5_571; w_5_572<=Wgt_5_572; w_5_573<=Wgt_5_573; w_5_574<=Wgt_5_574; w_5_575<=Wgt_5_575; w_5_576<=Wgt_5_576; w_5_577<=Wgt_5_577; w_5_578<=Wgt_5_578; w_5_579<=Wgt_5_579; w_5_580<=Wgt_5_580; w_5_581<=Wgt_5_581; w_5_582<=Wgt_5_582; w_5_583<=Wgt_5_583; w_5_584<=Wgt_5_584; w_5_585<=Wgt_5_585; w_5_586<=Wgt_5_586; w_5_587<=Wgt_5_587; w_5_588<=Wgt_5_588; w_5_589<=Wgt_5_589; w_5_590<=Wgt_5_590; w_5_591<=Wgt_5_591; w_5_592<=Wgt_5_592; w_5_593<=Wgt_5_593; w_5_594<=Wgt_5_594; w_5_595<=Wgt_5_595; w_5_596<=Wgt_5_596; w_5_597<=Wgt_5_597; w_5_598<=Wgt_5_598; w_5_599<=Wgt_5_599; w_5_600<=Wgt_5_600; w_5_601<=Wgt_5_601; w_5_602<=Wgt_5_602; w_5_603<=Wgt_5_603; w_5_604<=Wgt_5_604; w_5_605<=Wgt_5_605; w_5_606<=Wgt_5_606; w_5_607<=Wgt_5_607; w_5_608<=Wgt_5_608; w_5_609<=Wgt_5_609; w_5_610<=Wgt_5_610; w_5_611<=Wgt_5_611; w_5_612<=Wgt_5_612; w_5_613<=Wgt_5_613; w_5_614<=Wgt_5_614; w_5_615<=Wgt_5_615; w_5_616<=Wgt_5_616; w_5_617<=Wgt_5_617; w_5_618<=Wgt_5_618; w_5_619<=Wgt_5_619; w_5_620<=Wgt_5_620; w_5_621<=Wgt_5_621; w_5_622<=Wgt_5_622; w_5_623<=Wgt_5_623; w_5_624<=Wgt_5_624; w_5_625<=Wgt_5_625; w_5_626<=Wgt_5_626; w_5_627<=Wgt_5_627; w_5_628<=Wgt_5_628; w_5_629<=Wgt_5_629; w_5_630<=Wgt_5_630; w_5_631<=Wgt_5_631; w_5_632<=Wgt_5_632; w_5_633<=Wgt_5_633; w_5_634<=Wgt_5_634; w_5_635<=Wgt_5_635; w_5_636<=Wgt_5_636; w_5_637<=Wgt_5_637; w_5_638<=Wgt_5_638; w_5_639<=Wgt_5_639; w_5_640<=Wgt_5_640; w_5_641<=Wgt_5_641; w_5_642<=Wgt_5_642; w_5_643<=Wgt_5_643; w_5_644<=Wgt_5_644; w_5_645<=Wgt_5_645; w_5_646<=Wgt_5_646; w_5_647<=Wgt_5_647; w_5_648<=Wgt_5_648; w_5_649<=Wgt_5_649; w_5_650<=Wgt_5_650; w_5_651<=Wgt_5_651; w_5_652<=Wgt_5_652; w_5_653<=Wgt_5_653; w_5_654<=Wgt_5_654; w_5_655<=Wgt_5_655; w_5_656<=Wgt_5_656; w_5_657<=Wgt_5_657; w_5_658<=Wgt_5_658; w_5_659<=Wgt_5_659; w_5_660<=Wgt_5_660; w_5_661<=Wgt_5_661; w_5_662<=Wgt_5_662; w_5_663<=Wgt_5_663; w_5_664<=Wgt_5_664; w_5_665<=Wgt_5_665; w_5_666<=Wgt_5_666; w_5_667<=Wgt_5_667; w_5_668<=Wgt_5_668; w_5_669<=Wgt_5_669; w_5_670<=Wgt_5_670; w_5_671<=Wgt_5_671; w_5_672<=Wgt_5_672; w_5_673<=Wgt_5_673; w_5_674<=Wgt_5_674; w_5_675<=Wgt_5_675; w_5_676<=Wgt_5_676; w_5_677<=Wgt_5_677; w_5_678<=Wgt_5_678; w_5_679<=Wgt_5_679; w_5_680<=Wgt_5_680; w_5_681<=Wgt_5_681; w_5_682<=Wgt_5_682; w_5_683<=Wgt_5_683; w_5_684<=Wgt_5_684; w_5_685<=Wgt_5_685; w_5_686<=Wgt_5_686; w_5_687<=Wgt_5_687; w_5_688<=Wgt_5_688; w_5_689<=Wgt_5_689; w_5_690<=Wgt_5_690; w_5_691<=Wgt_5_691; w_5_692<=Wgt_5_692; w_5_693<=Wgt_5_693; w_5_694<=Wgt_5_694; w_5_695<=Wgt_5_695; w_5_696<=Wgt_5_696; w_5_697<=Wgt_5_697; w_5_698<=Wgt_5_698; w_5_699<=Wgt_5_699; w_5_700<=Wgt_5_700; w_5_701<=Wgt_5_701; w_5_702<=Wgt_5_702; w_5_703<=Wgt_5_703; w_5_704<=Wgt_5_704; w_5_705<=Wgt_5_705; w_5_706<=Wgt_5_706; w_5_707<=Wgt_5_707; w_5_708<=Wgt_5_708; w_5_709<=Wgt_5_709; w_5_710<=Wgt_5_710; w_5_711<=Wgt_5_711; w_5_712<=Wgt_5_712; w_5_713<=Wgt_5_713; w_5_714<=Wgt_5_714; w_5_715<=Wgt_5_715; w_5_716<=Wgt_5_716; w_5_717<=Wgt_5_717; w_5_718<=Wgt_5_718; w_5_719<=Wgt_5_719; w_5_720<=Wgt_5_720; w_5_721<=Wgt_5_721; w_5_722<=Wgt_5_722; w_5_723<=Wgt_5_723; w_5_724<=Wgt_5_724; w_5_725<=Wgt_5_725; w_5_726<=Wgt_5_726; w_5_727<=Wgt_5_727; w_5_728<=Wgt_5_728; w_5_729<=Wgt_5_729; w_5_730<=Wgt_5_730; w_5_731<=Wgt_5_731; w_5_732<=Wgt_5_732; w_5_733<=Wgt_5_733; w_5_734<=Wgt_5_734; w_5_735<=Wgt_5_735; w_5_736<=Wgt_5_736; w_5_737<=Wgt_5_737; w_5_738<=Wgt_5_738; w_5_739<=Wgt_5_739; w_5_740<=Wgt_5_740; w_5_741<=Wgt_5_741; w_5_742<=Wgt_5_742; w_5_743<=Wgt_5_743; w_5_744<=Wgt_5_744; w_5_745<=Wgt_5_745; w_5_746<=Wgt_5_746; w_5_747<=Wgt_5_747; w_5_748<=Wgt_5_748; w_5_749<=Wgt_5_749; w_5_750<=Wgt_5_750; w_5_751<=Wgt_5_751; w_5_752<=Wgt_5_752; w_5_753<=Wgt_5_753; w_5_754<=Wgt_5_754; w_5_755<=Wgt_5_755; w_5_756<=Wgt_5_756; w_5_757<=Wgt_5_757; w_5_758<=Wgt_5_758; w_5_759<=Wgt_5_759; w_5_760<=Wgt_5_760; w_5_761<=Wgt_5_761; w_5_762<=Wgt_5_762; w_5_763<=Wgt_5_763; w_5_764<=Wgt_5_764; w_5_765<=Wgt_5_765; w_5_766<=Wgt_5_766; w_5_767<=Wgt_5_767; w_5_768<=Wgt_5_768; w_5_769<=Wgt_5_769; w_5_770<=Wgt_5_770; w_5_771<=Wgt_5_771; w_5_772<=Wgt_5_772; w_5_773<=Wgt_5_773; w_5_774<=Wgt_5_774; w_5_775<=Wgt_5_775; w_5_776<=Wgt_5_776; w_5_777<=Wgt_5_777; w_5_778<=Wgt_5_778; w_5_779<=Wgt_5_779; w_5_780<=Wgt_5_780; w_5_781<=Wgt_5_781; w_5_782<=Wgt_5_782; w_5_783<=Wgt_5_783; w_5_784<=Wgt_5_784; 
					w_6_0<=Wgt_6_0; w_6_1<=Wgt_6_1; w_6_2<=Wgt_6_2; w_6_3<=Wgt_6_3; w_6_4<=Wgt_6_4; w_6_5<=Wgt_6_5; w_6_6<=Wgt_6_6; w_6_7<=Wgt_6_7; w_6_8<=Wgt_6_8; w_6_9<=Wgt_6_9; w_6_10<=Wgt_6_10; w_6_11<=Wgt_6_11; w_6_12<=Wgt_6_12; w_6_13<=Wgt_6_13; w_6_14<=Wgt_6_14; w_6_15<=Wgt_6_15; w_6_16<=Wgt_6_16; w_6_17<=Wgt_6_17; w_6_18<=Wgt_6_18; w_6_19<=Wgt_6_19; w_6_20<=Wgt_6_20; w_6_21<=Wgt_6_21; w_6_22<=Wgt_6_22; w_6_23<=Wgt_6_23; w_6_24<=Wgt_6_24; w_6_25<=Wgt_6_25; w_6_26<=Wgt_6_26; w_6_27<=Wgt_6_27; w_6_28<=Wgt_6_28; w_6_29<=Wgt_6_29; w_6_30<=Wgt_6_30; w_6_31<=Wgt_6_31; w_6_32<=Wgt_6_32; w_6_33<=Wgt_6_33; w_6_34<=Wgt_6_34; w_6_35<=Wgt_6_35; w_6_36<=Wgt_6_36; w_6_37<=Wgt_6_37; w_6_38<=Wgt_6_38; w_6_39<=Wgt_6_39; w_6_40<=Wgt_6_40; w_6_41<=Wgt_6_41; w_6_42<=Wgt_6_42; w_6_43<=Wgt_6_43; w_6_44<=Wgt_6_44; w_6_45<=Wgt_6_45; w_6_46<=Wgt_6_46; w_6_47<=Wgt_6_47; w_6_48<=Wgt_6_48; w_6_49<=Wgt_6_49; w_6_50<=Wgt_6_50; w_6_51<=Wgt_6_51; w_6_52<=Wgt_6_52; w_6_53<=Wgt_6_53; w_6_54<=Wgt_6_54; w_6_55<=Wgt_6_55; w_6_56<=Wgt_6_56; w_6_57<=Wgt_6_57; w_6_58<=Wgt_6_58; w_6_59<=Wgt_6_59; w_6_60<=Wgt_6_60; w_6_61<=Wgt_6_61; w_6_62<=Wgt_6_62; w_6_63<=Wgt_6_63; w_6_64<=Wgt_6_64; w_6_65<=Wgt_6_65; w_6_66<=Wgt_6_66; w_6_67<=Wgt_6_67; w_6_68<=Wgt_6_68; w_6_69<=Wgt_6_69; w_6_70<=Wgt_6_70; w_6_71<=Wgt_6_71; w_6_72<=Wgt_6_72; w_6_73<=Wgt_6_73; w_6_74<=Wgt_6_74; w_6_75<=Wgt_6_75; w_6_76<=Wgt_6_76; w_6_77<=Wgt_6_77; w_6_78<=Wgt_6_78; w_6_79<=Wgt_6_79; w_6_80<=Wgt_6_80; w_6_81<=Wgt_6_81; w_6_82<=Wgt_6_82; w_6_83<=Wgt_6_83; w_6_84<=Wgt_6_84; w_6_85<=Wgt_6_85; w_6_86<=Wgt_6_86; w_6_87<=Wgt_6_87; w_6_88<=Wgt_6_88; w_6_89<=Wgt_6_89; w_6_90<=Wgt_6_90; w_6_91<=Wgt_6_91; w_6_92<=Wgt_6_92; w_6_93<=Wgt_6_93; w_6_94<=Wgt_6_94; w_6_95<=Wgt_6_95; w_6_96<=Wgt_6_96; w_6_97<=Wgt_6_97; w_6_98<=Wgt_6_98; w_6_99<=Wgt_6_99; w_6_100<=Wgt_6_100; w_6_101<=Wgt_6_101; w_6_102<=Wgt_6_102; w_6_103<=Wgt_6_103; w_6_104<=Wgt_6_104; w_6_105<=Wgt_6_105; w_6_106<=Wgt_6_106; w_6_107<=Wgt_6_107; w_6_108<=Wgt_6_108; w_6_109<=Wgt_6_109; w_6_110<=Wgt_6_110; w_6_111<=Wgt_6_111; w_6_112<=Wgt_6_112; w_6_113<=Wgt_6_113; w_6_114<=Wgt_6_114; w_6_115<=Wgt_6_115; w_6_116<=Wgt_6_116; w_6_117<=Wgt_6_117; w_6_118<=Wgt_6_118; w_6_119<=Wgt_6_119; w_6_120<=Wgt_6_120; w_6_121<=Wgt_6_121; w_6_122<=Wgt_6_122; w_6_123<=Wgt_6_123; w_6_124<=Wgt_6_124; w_6_125<=Wgt_6_125; w_6_126<=Wgt_6_126; w_6_127<=Wgt_6_127; w_6_128<=Wgt_6_128; w_6_129<=Wgt_6_129; w_6_130<=Wgt_6_130; w_6_131<=Wgt_6_131; w_6_132<=Wgt_6_132; w_6_133<=Wgt_6_133; w_6_134<=Wgt_6_134; w_6_135<=Wgt_6_135; w_6_136<=Wgt_6_136; w_6_137<=Wgt_6_137; w_6_138<=Wgt_6_138; w_6_139<=Wgt_6_139; w_6_140<=Wgt_6_140; w_6_141<=Wgt_6_141; w_6_142<=Wgt_6_142; w_6_143<=Wgt_6_143; w_6_144<=Wgt_6_144; w_6_145<=Wgt_6_145; w_6_146<=Wgt_6_146; w_6_147<=Wgt_6_147; w_6_148<=Wgt_6_148; w_6_149<=Wgt_6_149; w_6_150<=Wgt_6_150; w_6_151<=Wgt_6_151; w_6_152<=Wgt_6_152; w_6_153<=Wgt_6_153; w_6_154<=Wgt_6_154; w_6_155<=Wgt_6_155; w_6_156<=Wgt_6_156; w_6_157<=Wgt_6_157; w_6_158<=Wgt_6_158; w_6_159<=Wgt_6_159; w_6_160<=Wgt_6_160; w_6_161<=Wgt_6_161; w_6_162<=Wgt_6_162; w_6_163<=Wgt_6_163; w_6_164<=Wgt_6_164; w_6_165<=Wgt_6_165; w_6_166<=Wgt_6_166; w_6_167<=Wgt_6_167; w_6_168<=Wgt_6_168; w_6_169<=Wgt_6_169; w_6_170<=Wgt_6_170; w_6_171<=Wgt_6_171; w_6_172<=Wgt_6_172; w_6_173<=Wgt_6_173; w_6_174<=Wgt_6_174; w_6_175<=Wgt_6_175; w_6_176<=Wgt_6_176; w_6_177<=Wgt_6_177; w_6_178<=Wgt_6_178; w_6_179<=Wgt_6_179; w_6_180<=Wgt_6_180; w_6_181<=Wgt_6_181; w_6_182<=Wgt_6_182; w_6_183<=Wgt_6_183; w_6_184<=Wgt_6_184; w_6_185<=Wgt_6_185; w_6_186<=Wgt_6_186; w_6_187<=Wgt_6_187; w_6_188<=Wgt_6_188; w_6_189<=Wgt_6_189; w_6_190<=Wgt_6_190; w_6_191<=Wgt_6_191; w_6_192<=Wgt_6_192; w_6_193<=Wgt_6_193; w_6_194<=Wgt_6_194; w_6_195<=Wgt_6_195; w_6_196<=Wgt_6_196; w_6_197<=Wgt_6_197; w_6_198<=Wgt_6_198; w_6_199<=Wgt_6_199; w_6_200<=Wgt_6_200; w_6_201<=Wgt_6_201; w_6_202<=Wgt_6_202; w_6_203<=Wgt_6_203; w_6_204<=Wgt_6_204; w_6_205<=Wgt_6_205; w_6_206<=Wgt_6_206; w_6_207<=Wgt_6_207; w_6_208<=Wgt_6_208; w_6_209<=Wgt_6_209; w_6_210<=Wgt_6_210; w_6_211<=Wgt_6_211; w_6_212<=Wgt_6_212; w_6_213<=Wgt_6_213; w_6_214<=Wgt_6_214; w_6_215<=Wgt_6_215; w_6_216<=Wgt_6_216; w_6_217<=Wgt_6_217; w_6_218<=Wgt_6_218; w_6_219<=Wgt_6_219; w_6_220<=Wgt_6_220; w_6_221<=Wgt_6_221; w_6_222<=Wgt_6_222; w_6_223<=Wgt_6_223; w_6_224<=Wgt_6_224; w_6_225<=Wgt_6_225; w_6_226<=Wgt_6_226; w_6_227<=Wgt_6_227; w_6_228<=Wgt_6_228; w_6_229<=Wgt_6_229; w_6_230<=Wgt_6_230; w_6_231<=Wgt_6_231; w_6_232<=Wgt_6_232; w_6_233<=Wgt_6_233; w_6_234<=Wgt_6_234; w_6_235<=Wgt_6_235; w_6_236<=Wgt_6_236; w_6_237<=Wgt_6_237; w_6_238<=Wgt_6_238; w_6_239<=Wgt_6_239; w_6_240<=Wgt_6_240; w_6_241<=Wgt_6_241; w_6_242<=Wgt_6_242; w_6_243<=Wgt_6_243; w_6_244<=Wgt_6_244; w_6_245<=Wgt_6_245; w_6_246<=Wgt_6_246; w_6_247<=Wgt_6_247; w_6_248<=Wgt_6_248; w_6_249<=Wgt_6_249; w_6_250<=Wgt_6_250; w_6_251<=Wgt_6_251; w_6_252<=Wgt_6_252; w_6_253<=Wgt_6_253; w_6_254<=Wgt_6_254; w_6_255<=Wgt_6_255; w_6_256<=Wgt_6_256; w_6_257<=Wgt_6_257; w_6_258<=Wgt_6_258; w_6_259<=Wgt_6_259; w_6_260<=Wgt_6_260; w_6_261<=Wgt_6_261; w_6_262<=Wgt_6_262; w_6_263<=Wgt_6_263; w_6_264<=Wgt_6_264; w_6_265<=Wgt_6_265; w_6_266<=Wgt_6_266; w_6_267<=Wgt_6_267; w_6_268<=Wgt_6_268; w_6_269<=Wgt_6_269; w_6_270<=Wgt_6_270; w_6_271<=Wgt_6_271; w_6_272<=Wgt_6_272; w_6_273<=Wgt_6_273; w_6_274<=Wgt_6_274; w_6_275<=Wgt_6_275; w_6_276<=Wgt_6_276; w_6_277<=Wgt_6_277; w_6_278<=Wgt_6_278; w_6_279<=Wgt_6_279; w_6_280<=Wgt_6_280; w_6_281<=Wgt_6_281; w_6_282<=Wgt_6_282; w_6_283<=Wgt_6_283; w_6_284<=Wgt_6_284; w_6_285<=Wgt_6_285; w_6_286<=Wgt_6_286; w_6_287<=Wgt_6_287; w_6_288<=Wgt_6_288; w_6_289<=Wgt_6_289; w_6_290<=Wgt_6_290; w_6_291<=Wgt_6_291; w_6_292<=Wgt_6_292; w_6_293<=Wgt_6_293; w_6_294<=Wgt_6_294; w_6_295<=Wgt_6_295; w_6_296<=Wgt_6_296; w_6_297<=Wgt_6_297; w_6_298<=Wgt_6_298; w_6_299<=Wgt_6_299; w_6_300<=Wgt_6_300; w_6_301<=Wgt_6_301; w_6_302<=Wgt_6_302; w_6_303<=Wgt_6_303; w_6_304<=Wgt_6_304; w_6_305<=Wgt_6_305; w_6_306<=Wgt_6_306; w_6_307<=Wgt_6_307; w_6_308<=Wgt_6_308; w_6_309<=Wgt_6_309; w_6_310<=Wgt_6_310; w_6_311<=Wgt_6_311; w_6_312<=Wgt_6_312; w_6_313<=Wgt_6_313; w_6_314<=Wgt_6_314; w_6_315<=Wgt_6_315; w_6_316<=Wgt_6_316; w_6_317<=Wgt_6_317; w_6_318<=Wgt_6_318; w_6_319<=Wgt_6_319; w_6_320<=Wgt_6_320; w_6_321<=Wgt_6_321; w_6_322<=Wgt_6_322; w_6_323<=Wgt_6_323; w_6_324<=Wgt_6_324; w_6_325<=Wgt_6_325; w_6_326<=Wgt_6_326; w_6_327<=Wgt_6_327; w_6_328<=Wgt_6_328; w_6_329<=Wgt_6_329; w_6_330<=Wgt_6_330; w_6_331<=Wgt_6_331; w_6_332<=Wgt_6_332; w_6_333<=Wgt_6_333; w_6_334<=Wgt_6_334; w_6_335<=Wgt_6_335; w_6_336<=Wgt_6_336; w_6_337<=Wgt_6_337; w_6_338<=Wgt_6_338; w_6_339<=Wgt_6_339; w_6_340<=Wgt_6_340; w_6_341<=Wgt_6_341; w_6_342<=Wgt_6_342; w_6_343<=Wgt_6_343; w_6_344<=Wgt_6_344; w_6_345<=Wgt_6_345; w_6_346<=Wgt_6_346; w_6_347<=Wgt_6_347; w_6_348<=Wgt_6_348; w_6_349<=Wgt_6_349; w_6_350<=Wgt_6_350; w_6_351<=Wgt_6_351; w_6_352<=Wgt_6_352; w_6_353<=Wgt_6_353; w_6_354<=Wgt_6_354; w_6_355<=Wgt_6_355; w_6_356<=Wgt_6_356; w_6_357<=Wgt_6_357; w_6_358<=Wgt_6_358; w_6_359<=Wgt_6_359; w_6_360<=Wgt_6_360; w_6_361<=Wgt_6_361; w_6_362<=Wgt_6_362; w_6_363<=Wgt_6_363; w_6_364<=Wgt_6_364; w_6_365<=Wgt_6_365; w_6_366<=Wgt_6_366; w_6_367<=Wgt_6_367; w_6_368<=Wgt_6_368; w_6_369<=Wgt_6_369; w_6_370<=Wgt_6_370; w_6_371<=Wgt_6_371; w_6_372<=Wgt_6_372; w_6_373<=Wgt_6_373; w_6_374<=Wgt_6_374; w_6_375<=Wgt_6_375; w_6_376<=Wgt_6_376; w_6_377<=Wgt_6_377; w_6_378<=Wgt_6_378; w_6_379<=Wgt_6_379; w_6_380<=Wgt_6_380; w_6_381<=Wgt_6_381; w_6_382<=Wgt_6_382; w_6_383<=Wgt_6_383; w_6_384<=Wgt_6_384; w_6_385<=Wgt_6_385; w_6_386<=Wgt_6_386; w_6_387<=Wgt_6_387; w_6_388<=Wgt_6_388; w_6_389<=Wgt_6_389; w_6_390<=Wgt_6_390; w_6_391<=Wgt_6_391; w_6_392<=Wgt_6_392; w_6_393<=Wgt_6_393; w_6_394<=Wgt_6_394; w_6_395<=Wgt_6_395; w_6_396<=Wgt_6_396; w_6_397<=Wgt_6_397; w_6_398<=Wgt_6_398; w_6_399<=Wgt_6_399; w_6_400<=Wgt_6_400; w_6_401<=Wgt_6_401; w_6_402<=Wgt_6_402; w_6_403<=Wgt_6_403; w_6_404<=Wgt_6_404; w_6_405<=Wgt_6_405; w_6_406<=Wgt_6_406; w_6_407<=Wgt_6_407; w_6_408<=Wgt_6_408; w_6_409<=Wgt_6_409; w_6_410<=Wgt_6_410; w_6_411<=Wgt_6_411; w_6_412<=Wgt_6_412; w_6_413<=Wgt_6_413; w_6_414<=Wgt_6_414; w_6_415<=Wgt_6_415; w_6_416<=Wgt_6_416; w_6_417<=Wgt_6_417; w_6_418<=Wgt_6_418; w_6_419<=Wgt_6_419; w_6_420<=Wgt_6_420; w_6_421<=Wgt_6_421; w_6_422<=Wgt_6_422; w_6_423<=Wgt_6_423; w_6_424<=Wgt_6_424; w_6_425<=Wgt_6_425; w_6_426<=Wgt_6_426; w_6_427<=Wgt_6_427; w_6_428<=Wgt_6_428; w_6_429<=Wgt_6_429; w_6_430<=Wgt_6_430; w_6_431<=Wgt_6_431; w_6_432<=Wgt_6_432; w_6_433<=Wgt_6_433; w_6_434<=Wgt_6_434; w_6_435<=Wgt_6_435; w_6_436<=Wgt_6_436; w_6_437<=Wgt_6_437; w_6_438<=Wgt_6_438; w_6_439<=Wgt_6_439; w_6_440<=Wgt_6_440; w_6_441<=Wgt_6_441; w_6_442<=Wgt_6_442; w_6_443<=Wgt_6_443; w_6_444<=Wgt_6_444; w_6_445<=Wgt_6_445; w_6_446<=Wgt_6_446; w_6_447<=Wgt_6_447; w_6_448<=Wgt_6_448; w_6_449<=Wgt_6_449; w_6_450<=Wgt_6_450; w_6_451<=Wgt_6_451; w_6_452<=Wgt_6_452; w_6_453<=Wgt_6_453; w_6_454<=Wgt_6_454; w_6_455<=Wgt_6_455; w_6_456<=Wgt_6_456; w_6_457<=Wgt_6_457; w_6_458<=Wgt_6_458; w_6_459<=Wgt_6_459; w_6_460<=Wgt_6_460; w_6_461<=Wgt_6_461; w_6_462<=Wgt_6_462; w_6_463<=Wgt_6_463; w_6_464<=Wgt_6_464; w_6_465<=Wgt_6_465; w_6_466<=Wgt_6_466; w_6_467<=Wgt_6_467; w_6_468<=Wgt_6_468; w_6_469<=Wgt_6_469; w_6_470<=Wgt_6_470; w_6_471<=Wgt_6_471; w_6_472<=Wgt_6_472; w_6_473<=Wgt_6_473; w_6_474<=Wgt_6_474; w_6_475<=Wgt_6_475; w_6_476<=Wgt_6_476; w_6_477<=Wgt_6_477; w_6_478<=Wgt_6_478; w_6_479<=Wgt_6_479; w_6_480<=Wgt_6_480; w_6_481<=Wgt_6_481; w_6_482<=Wgt_6_482; w_6_483<=Wgt_6_483; w_6_484<=Wgt_6_484; w_6_485<=Wgt_6_485; w_6_486<=Wgt_6_486; w_6_487<=Wgt_6_487; w_6_488<=Wgt_6_488; w_6_489<=Wgt_6_489; w_6_490<=Wgt_6_490; w_6_491<=Wgt_6_491; w_6_492<=Wgt_6_492; w_6_493<=Wgt_6_493; w_6_494<=Wgt_6_494; w_6_495<=Wgt_6_495; w_6_496<=Wgt_6_496; w_6_497<=Wgt_6_497; w_6_498<=Wgt_6_498; w_6_499<=Wgt_6_499; w_6_500<=Wgt_6_500; w_6_501<=Wgt_6_501; w_6_502<=Wgt_6_502; w_6_503<=Wgt_6_503; w_6_504<=Wgt_6_504; w_6_505<=Wgt_6_505; w_6_506<=Wgt_6_506; w_6_507<=Wgt_6_507; w_6_508<=Wgt_6_508; w_6_509<=Wgt_6_509; w_6_510<=Wgt_6_510; w_6_511<=Wgt_6_511; w_6_512<=Wgt_6_512; w_6_513<=Wgt_6_513; w_6_514<=Wgt_6_514; w_6_515<=Wgt_6_515; w_6_516<=Wgt_6_516; w_6_517<=Wgt_6_517; w_6_518<=Wgt_6_518; w_6_519<=Wgt_6_519; w_6_520<=Wgt_6_520; w_6_521<=Wgt_6_521; w_6_522<=Wgt_6_522; w_6_523<=Wgt_6_523; w_6_524<=Wgt_6_524; w_6_525<=Wgt_6_525; w_6_526<=Wgt_6_526; w_6_527<=Wgt_6_527; w_6_528<=Wgt_6_528; w_6_529<=Wgt_6_529; w_6_530<=Wgt_6_530; w_6_531<=Wgt_6_531; w_6_532<=Wgt_6_532; w_6_533<=Wgt_6_533; w_6_534<=Wgt_6_534; w_6_535<=Wgt_6_535; w_6_536<=Wgt_6_536; w_6_537<=Wgt_6_537; w_6_538<=Wgt_6_538; w_6_539<=Wgt_6_539; w_6_540<=Wgt_6_540; w_6_541<=Wgt_6_541; w_6_542<=Wgt_6_542; w_6_543<=Wgt_6_543; w_6_544<=Wgt_6_544; w_6_545<=Wgt_6_545; w_6_546<=Wgt_6_546; w_6_547<=Wgt_6_547; w_6_548<=Wgt_6_548; w_6_549<=Wgt_6_549; w_6_550<=Wgt_6_550; w_6_551<=Wgt_6_551; w_6_552<=Wgt_6_552; w_6_553<=Wgt_6_553; w_6_554<=Wgt_6_554; w_6_555<=Wgt_6_555; w_6_556<=Wgt_6_556; w_6_557<=Wgt_6_557; w_6_558<=Wgt_6_558; w_6_559<=Wgt_6_559; w_6_560<=Wgt_6_560; w_6_561<=Wgt_6_561; w_6_562<=Wgt_6_562; w_6_563<=Wgt_6_563; w_6_564<=Wgt_6_564; w_6_565<=Wgt_6_565; w_6_566<=Wgt_6_566; w_6_567<=Wgt_6_567; w_6_568<=Wgt_6_568; w_6_569<=Wgt_6_569; w_6_570<=Wgt_6_570; w_6_571<=Wgt_6_571; w_6_572<=Wgt_6_572; w_6_573<=Wgt_6_573; w_6_574<=Wgt_6_574; w_6_575<=Wgt_6_575; w_6_576<=Wgt_6_576; w_6_577<=Wgt_6_577; w_6_578<=Wgt_6_578; w_6_579<=Wgt_6_579; w_6_580<=Wgt_6_580; w_6_581<=Wgt_6_581; w_6_582<=Wgt_6_582; w_6_583<=Wgt_6_583; w_6_584<=Wgt_6_584; w_6_585<=Wgt_6_585; w_6_586<=Wgt_6_586; w_6_587<=Wgt_6_587; w_6_588<=Wgt_6_588; w_6_589<=Wgt_6_589; w_6_590<=Wgt_6_590; w_6_591<=Wgt_6_591; w_6_592<=Wgt_6_592; w_6_593<=Wgt_6_593; w_6_594<=Wgt_6_594; w_6_595<=Wgt_6_595; w_6_596<=Wgt_6_596; w_6_597<=Wgt_6_597; w_6_598<=Wgt_6_598; w_6_599<=Wgt_6_599; w_6_600<=Wgt_6_600; w_6_601<=Wgt_6_601; w_6_602<=Wgt_6_602; w_6_603<=Wgt_6_603; w_6_604<=Wgt_6_604; w_6_605<=Wgt_6_605; w_6_606<=Wgt_6_606; w_6_607<=Wgt_6_607; w_6_608<=Wgt_6_608; w_6_609<=Wgt_6_609; w_6_610<=Wgt_6_610; w_6_611<=Wgt_6_611; w_6_612<=Wgt_6_612; w_6_613<=Wgt_6_613; w_6_614<=Wgt_6_614; w_6_615<=Wgt_6_615; w_6_616<=Wgt_6_616; w_6_617<=Wgt_6_617; w_6_618<=Wgt_6_618; w_6_619<=Wgt_6_619; w_6_620<=Wgt_6_620; w_6_621<=Wgt_6_621; w_6_622<=Wgt_6_622; w_6_623<=Wgt_6_623; w_6_624<=Wgt_6_624; w_6_625<=Wgt_6_625; w_6_626<=Wgt_6_626; w_6_627<=Wgt_6_627; w_6_628<=Wgt_6_628; w_6_629<=Wgt_6_629; w_6_630<=Wgt_6_630; w_6_631<=Wgt_6_631; w_6_632<=Wgt_6_632; w_6_633<=Wgt_6_633; w_6_634<=Wgt_6_634; w_6_635<=Wgt_6_635; w_6_636<=Wgt_6_636; w_6_637<=Wgt_6_637; w_6_638<=Wgt_6_638; w_6_639<=Wgt_6_639; w_6_640<=Wgt_6_640; w_6_641<=Wgt_6_641; w_6_642<=Wgt_6_642; w_6_643<=Wgt_6_643; w_6_644<=Wgt_6_644; w_6_645<=Wgt_6_645; w_6_646<=Wgt_6_646; w_6_647<=Wgt_6_647; w_6_648<=Wgt_6_648; w_6_649<=Wgt_6_649; w_6_650<=Wgt_6_650; w_6_651<=Wgt_6_651; w_6_652<=Wgt_6_652; w_6_653<=Wgt_6_653; w_6_654<=Wgt_6_654; w_6_655<=Wgt_6_655; w_6_656<=Wgt_6_656; w_6_657<=Wgt_6_657; w_6_658<=Wgt_6_658; w_6_659<=Wgt_6_659; w_6_660<=Wgt_6_660; w_6_661<=Wgt_6_661; w_6_662<=Wgt_6_662; w_6_663<=Wgt_6_663; w_6_664<=Wgt_6_664; w_6_665<=Wgt_6_665; w_6_666<=Wgt_6_666; w_6_667<=Wgt_6_667; w_6_668<=Wgt_6_668; w_6_669<=Wgt_6_669; w_6_670<=Wgt_6_670; w_6_671<=Wgt_6_671; w_6_672<=Wgt_6_672; w_6_673<=Wgt_6_673; w_6_674<=Wgt_6_674; w_6_675<=Wgt_6_675; w_6_676<=Wgt_6_676; w_6_677<=Wgt_6_677; w_6_678<=Wgt_6_678; w_6_679<=Wgt_6_679; w_6_680<=Wgt_6_680; w_6_681<=Wgt_6_681; w_6_682<=Wgt_6_682; w_6_683<=Wgt_6_683; w_6_684<=Wgt_6_684; w_6_685<=Wgt_6_685; w_6_686<=Wgt_6_686; w_6_687<=Wgt_6_687; w_6_688<=Wgt_6_688; w_6_689<=Wgt_6_689; w_6_690<=Wgt_6_690; w_6_691<=Wgt_6_691; w_6_692<=Wgt_6_692; w_6_693<=Wgt_6_693; w_6_694<=Wgt_6_694; w_6_695<=Wgt_6_695; w_6_696<=Wgt_6_696; w_6_697<=Wgt_6_697; w_6_698<=Wgt_6_698; w_6_699<=Wgt_6_699; w_6_700<=Wgt_6_700; w_6_701<=Wgt_6_701; w_6_702<=Wgt_6_702; w_6_703<=Wgt_6_703; w_6_704<=Wgt_6_704; w_6_705<=Wgt_6_705; w_6_706<=Wgt_6_706; w_6_707<=Wgt_6_707; w_6_708<=Wgt_6_708; w_6_709<=Wgt_6_709; w_6_710<=Wgt_6_710; w_6_711<=Wgt_6_711; w_6_712<=Wgt_6_712; w_6_713<=Wgt_6_713; w_6_714<=Wgt_6_714; w_6_715<=Wgt_6_715; w_6_716<=Wgt_6_716; w_6_717<=Wgt_6_717; w_6_718<=Wgt_6_718; w_6_719<=Wgt_6_719; w_6_720<=Wgt_6_720; w_6_721<=Wgt_6_721; w_6_722<=Wgt_6_722; w_6_723<=Wgt_6_723; w_6_724<=Wgt_6_724; w_6_725<=Wgt_6_725; w_6_726<=Wgt_6_726; w_6_727<=Wgt_6_727; w_6_728<=Wgt_6_728; w_6_729<=Wgt_6_729; w_6_730<=Wgt_6_730; w_6_731<=Wgt_6_731; w_6_732<=Wgt_6_732; w_6_733<=Wgt_6_733; w_6_734<=Wgt_6_734; w_6_735<=Wgt_6_735; w_6_736<=Wgt_6_736; w_6_737<=Wgt_6_737; w_6_738<=Wgt_6_738; w_6_739<=Wgt_6_739; w_6_740<=Wgt_6_740; w_6_741<=Wgt_6_741; w_6_742<=Wgt_6_742; w_6_743<=Wgt_6_743; w_6_744<=Wgt_6_744; w_6_745<=Wgt_6_745; w_6_746<=Wgt_6_746; w_6_747<=Wgt_6_747; w_6_748<=Wgt_6_748; w_6_749<=Wgt_6_749; w_6_750<=Wgt_6_750; w_6_751<=Wgt_6_751; w_6_752<=Wgt_6_752; w_6_753<=Wgt_6_753; w_6_754<=Wgt_6_754; w_6_755<=Wgt_6_755; w_6_756<=Wgt_6_756; w_6_757<=Wgt_6_757; w_6_758<=Wgt_6_758; w_6_759<=Wgt_6_759; w_6_760<=Wgt_6_760; w_6_761<=Wgt_6_761; w_6_762<=Wgt_6_762; w_6_763<=Wgt_6_763; w_6_764<=Wgt_6_764; w_6_765<=Wgt_6_765; w_6_766<=Wgt_6_766; w_6_767<=Wgt_6_767; w_6_768<=Wgt_6_768; w_6_769<=Wgt_6_769; w_6_770<=Wgt_6_770; w_6_771<=Wgt_6_771; w_6_772<=Wgt_6_772; w_6_773<=Wgt_6_773; w_6_774<=Wgt_6_774; w_6_775<=Wgt_6_775; w_6_776<=Wgt_6_776; w_6_777<=Wgt_6_777; w_6_778<=Wgt_6_778; w_6_779<=Wgt_6_779; w_6_780<=Wgt_6_780; w_6_781<=Wgt_6_781; w_6_782<=Wgt_6_782; w_6_783<=Wgt_6_783; w_6_784<=Wgt_6_784; 
					w_7_0<=Wgt_7_0; w_7_1<=Wgt_7_1; w_7_2<=Wgt_7_2; w_7_3<=Wgt_7_3; w_7_4<=Wgt_7_4; w_7_5<=Wgt_7_5; w_7_6<=Wgt_7_6; w_7_7<=Wgt_7_7; w_7_8<=Wgt_7_8; w_7_9<=Wgt_7_9; w_7_10<=Wgt_7_10; w_7_11<=Wgt_7_11; w_7_12<=Wgt_7_12; w_7_13<=Wgt_7_13; w_7_14<=Wgt_7_14; w_7_15<=Wgt_7_15; w_7_16<=Wgt_7_16; w_7_17<=Wgt_7_17; w_7_18<=Wgt_7_18; w_7_19<=Wgt_7_19; w_7_20<=Wgt_7_20; w_7_21<=Wgt_7_21; w_7_22<=Wgt_7_22; w_7_23<=Wgt_7_23; w_7_24<=Wgt_7_24; w_7_25<=Wgt_7_25; w_7_26<=Wgt_7_26; w_7_27<=Wgt_7_27; w_7_28<=Wgt_7_28; w_7_29<=Wgt_7_29; w_7_30<=Wgt_7_30; w_7_31<=Wgt_7_31; w_7_32<=Wgt_7_32; w_7_33<=Wgt_7_33; w_7_34<=Wgt_7_34; w_7_35<=Wgt_7_35; w_7_36<=Wgt_7_36; w_7_37<=Wgt_7_37; w_7_38<=Wgt_7_38; w_7_39<=Wgt_7_39; w_7_40<=Wgt_7_40; w_7_41<=Wgt_7_41; w_7_42<=Wgt_7_42; w_7_43<=Wgt_7_43; w_7_44<=Wgt_7_44; w_7_45<=Wgt_7_45; w_7_46<=Wgt_7_46; w_7_47<=Wgt_7_47; w_7_48<=Wgt_7_48; w_7_49<=Wgt_7_49; w_7_50<=Wgt_7_50; w_7_51<=Wgt_7_51; w_7_52<=Wgt_7_52; w_7_53<=Wgt_7_53; w_7_54<=Wgt_7_54; w_7_55<=Wgt_7_55; w_7_56<=Wgt_7_56; w_7_57<=Wgt_7_57; w_7_58<=Wgt_7_58; w_7_59<=Wgt_7_59; w_7_60<=Wgt_7_60; w_7_61<=Wgt_7_61; w_7_62<=Wgt_7_62; w_7_63<=Wgt_7_63; w_7_64<=Wgt_7_64; w_7_65<=Wgt_7_65; w_7_66<=Wgt_7_66; w_7_67<=Wgt_7_67; w_7_68<=Wgt_7_68; w_7_69<=Wgt_7_69; w_7_70<=Wgt_7_70; w_7_71<=Wgt_7_71; w_7_72<=Wgt_7_72; w_7_73<=Wgt_7_73; w_7_74<=Wgt_7_74; w_7_75<=Wgt_7_75; w_7_76<=Wgt_7_76; w_7_77<=Wgt_7_77; w_7_78<=Wgt_7_78; w_7_79<=Wgt_7_79; w_7_80<=Wgt_7_80; w_7_81<=Wgt_7_81; w_7_82<=Wgt_7_82; w_7_83<=Wgt_7_83; w_7_84<=Wgt_7_84; w_7_85<=Wgt_7_85; w_7_86<=Wgt_7_86; w_7_87<=Wgt_7_87; w_7_88<=Wgt_7_88; w_7_89<=Wgt_7_89; w_7_90<=Wgt_7_90; w_7_91<=Wgt_7_91; w_7_92<=Wgt_7_92; w_7_93<=Wgt_7_93; w_7_94<=Wgt_7_94; w_7_95<=Wgt_7_95; w_7_96<=Wgt_7_96; w_7_97<=Wgt_7_97; w_7_98<=Wgt_7_98; w_7_99<=Wgt_7_99; w_7_100<=Wgt_7_100; w_7_101<=Wgt_7_101; w_7_102<=Wgt_7_102; w_7_103<=Wgt_7_103; w_7_104<=Wgt_7_104; w_7_105<=Wgt_7_105; w_7_106<=Wgt_7_106; w_7_107<=Wgt_7_107; w_7_108<=Wgt_7_108; w_7_109<=Wgt_7_109; w_7_110<=Wgt_7_110; w_7_111<=Wgt_7_111; w_7_112<=Wgt_7_112; w_7_113<=Wgt_7_113; w_7_114<=Wgt_7_114; w_7_115<=Wgt_7_115; w_7_116<=Wgt_7_116; w_7_117<=Wgt_7_117; w_7_118<=Wgt_7_118; w_7_119<=Wgt_7_119; w_7_120<=Wgt_7_120; w_7_121<=Wgt_7_121; w_7_122<=Wgt_7_122; w_7_123<=Wgt_7_123; w_7_124<=Wgt_7_124; w_7_125<=Wgt_7_125; w_7_126<=Wgt_7_126; w_7_127<=Wgt_7_127; w_7_128<=Wgt_7_128; w_7_129<=Wgt_7_129; w_7_130<=Wgt_7_130; w_7_131<=Wgt_7_131; w_7_132<=Wgt_7_132; w_7_133<=Wgt_7_133; w_7_134<=Wgt_7_134; w_7_135<=Wgt_7_135; w_7_136<=Wgt_7_136; w_7_137<=Wgt_7_137; w_7_138<=Wgt_7_138; w_7_139<=Wgt_7_139; w_7_140<=Wgt_7_140; w_7_141<=Wgt_7_141; w_7_142<=Wgt_7_142; w_7_143<=Wgt_7_143; w_7_144<=Wgt_7_144; w_7_145<=Wgt_7_145; w_7_146<=Wgt_7_146; w_7_147<=Wgt_7_147; w_7_148<=Wgt_7_148; w_7_149<=Wgt_7_149; w_7_150<=Wgt_7_150; w_7_151<=Wgt_7_151; w_7_152<=Wgt_7_152; w_7_153<=Wgt_7_153; w_7_154<=Wgt_7_154; w_7_155<=Wgt_7_155; w_7_156<=Wgt_7_156; w_7_157<=Wgt_7_157; w_7_158<=Wgt_7_158; w_7_159<=Wgt_7_159; w_7_160<=Wgt_7_160; w_7_161<=Wgt_7_161; w_7_162<=Wgt_7_162; w_7_163<=Wgt_7_163; w_7_164<=Wgt_7_164; w_7_165<=Wgt_7_165; w_7_166<=Wgt_7_166; w_7_167<=Wgt_7_167; w_7_168<=Wgt_7_168; w_7_169<=Wgt_7_169; w_7_170<=Wgt_7_170; w_7_171<=Wgt_7_171; w_7_172<=Wgt_7_172; w_7_173<=Wgt_7_173; w_7_174<=Wgt_7_174; w_7_175<=Wgt_7_175; w_7_176<=Wgt_7_176; w_7_177<=Wgt_7_177; w_7_178<=Wgt_7_178; w_7_179<=Wgt_7_179; w_7_180<=Wgt_7_180; w_7_181<=Wgt_7_181; w_7_182<=Wgt_7_182; w_7_183<=Wgt_7_183; w_7_184<=Wgt_7_184; w_7_185<=Wgt_7_185; w_7_186<=Wgt_7_186; w_7_187<=Wgt_7_187; w_7_188<=Wgt_7_188; w_7_189<=Wgt_7_189; w_7_190<=Wgt_7_190; w_7_191<=Wgt_7_191; w_7_192<=Wgt_7_192; w_7_193<=Wgt_7_193; w_7_194<=Wgt_7_194; w_7_195<=Wgt_7_195; w_7_196<=Wgt_7_196; w_7_197<=Wgt_7_197; w_7_198<=Wgt_7_198; w_7_199<=Wgt_7_199; w_7_200<=Wgt_7_200; w_7_201<=Wgt_7_201; w_7_202<=Wgt_7_202; w_7_203<=Wgt_7_203; w_7_204<=Wgt_7_204; w_7_205<=Wgt_7_205; w_7_206<=Wgt_7_206; w_7_207<=Wgt_7_207; w_7_208<=Wgt_7_208; w_7_209<=Wgt_7_209; w_7_210<=Wgt_7_210; w_7_211<=Wgt_7_211; w_7_212<=Wgt_7_212; w_7_213<=Wgt_7_213; w_7_214<=Wgt_7_214; w_7_215<=Wgt_7_215; w_7_216<=Wgt_7_216; w_7_217<=Wgt_7_217; w_7_218<=Wgt_7_218; w_7_219<=Wgt_7_219; w_7_220<=Wgt_7_220; w_7_221<=Wgt_7_221; w_7_222<=Wgt_7_222; w_7_223<=Wgt_7_223; w_7_224<=Wgt_7_224; w_7_225<=Wgt_7_225; w_7_226<=Wgt_7_226; w_7_227<=Wgt_7_227; w_7_228<=Wgt_7_228; w_7_229<=Wgt_7_229; w_7_230<=Wgt_7_230; w_7_231<=Wgt_7_231; w_7_232<=Wgt_7_232; w_7_233<=Wgt_7_233; w_7_234<=Wgt_7_234; w_7_235<=Wgt_7_235; w_7_236<=Wgt_7_236; w_7_237<=Wgt_7_237; w_7_238<=Wgt_7_238; w_7_239<=Wgt_7_239; w_7_240<=Wgt_7_240; w_7_241<=Wgt_7_241; w_7_242<=Wgt_7_242; w_7_243<=Wgt_7_243; w_7_244<=Wgt_7_244; w_7_245<=Wgt_7_245; w_7_246<=Wgt_7_246; w_7_247<=Wgt_7_247; w_7_248<=Wgt_7_248; w_7_249<=Wgt_7_249; w_7_250<=Wgt_7_250; w_7_251<=Wgt_7_251; w_7_252<=Wgt_7_252; w_7_253<=Wgt_7_253; w_7_254<=Wgt_7_254; w_7_255<=Wgt_7_255; w_7_256<=Wgt_7_256; w_7_257<=Wgt_7_257; w_7_258<=Wgt_7_258; w_7_259<=Wgt_7_259; w_7_260<=Wgt_7_260; w_7_261<=Wgt_7_261; w_7_262<=Wgt_7_262; w_7_263<=Wgt_7_263; w_7_264<=Wgt_7_264; w_7_265<=Wgt_7_265; w_7_266<=Wgt_7_266; w_7_267<=Wgt_7_267; w_7_268<=Wgt_7_268; w_7_269<=Wgt_7_269; w_7_270<=Wgt_7_270; w_7_271<=Wgt_7_271; w_7_272<=Wgt_7_272; w_7_273<=Wgt_7_273; w_7_274<=Wgt_7_274; w_7_275<=Wgt_7_275; w_7_276<=Wgt_7_276; w_7_277<=Wgt_7_277; w_7_278<=Wgt_7_278; w_7_279<=Wgt_7_279; w_7_280<=Wgt_7_280; w_7_281<=Wgt_7_281; w_7_282<=Wgt_7_282; w_7_283<=Wgt_7_283; w_7_284<=Wgt_7_284; w_7_285<=Wgt_7_285; w_7_286<=Wgt_7_286; w_7_287<=Wgt_7_287; w_7_288<=Wgt_7_288; w_7_289<=Wgt_7_289; w_7_290<=Wgt_7_290; w_7_291<=Wgt_7_291; w_7_292<=Wgt_7_292; w_7_293<=Wgt_7_293; w_7_294<=Wgt_7_294; w_7_295<=Wgt_7_295; w_7_296<=Wgt_7_296; w_7_297<=Wgt_7_297; w_7_298<=Wgt_7_298; w_7_299<=Wgt_7_299; w_7_300<=Wgt_7_300; w_7_301<=Wgt_7_301; w_7_302<=Wgt_7_302; w_7_303<=Wgt_7_303; w_7_304<=Wgt_7_304; w_7_305<=Wgt_7_305; w_7_306<=Wgt_7_306; w_7_307<=Wgt_7_307; w_7_308<=Wgt_7_308; w_7_309<=Wgt_7_309; w_7_310<=Wgt_7_310; w_7_311<=Wgt_7_311; w_7_312<=Wgt_7_312; w_7_313<=Wgt_7_313; w_7_314<=Wgt_7_314; w_7_315<=Wgt_7_315; w_7_316<=Wgt_7_316; w_7_317<=Wgt_7_317; w_7_318<=Wgt_7_318; w_7_319<=Wgt_7_319; w_7_320<=Wgt_7_320; w_7_321<=Wgt_7_321; w_7_322<=Wgt_7_322; w_7_323<=Wgt_7_323; w_7_324<=Wgt_7_324; w_7_325<=Wgt_7_325; w_7_326<=Wgt_7_326; w_7_327<=Wgt_7_327; w_7_328<=Wgt_7_328; w_7_329<=Wgt_7_329; w_7_330<=Wgt_7_330; w_7_331<=Wgt_7_331; w_7_332<=Wgt_7_332; w_7_333<=Wgt_7_333; w_7_334<=Wgt_7_334; w_7_335<=Wgt_7_335; w_7_336<=Wgt_7_336; w_7_337<=Wgt_7_337; w_7_338<=Wgt_7_338; w_7_339<=Wgt_7_339; w_7_340<=Wgt_7_340; w_7_341<=Wgt_7_341; w_7_342<=Wgt_7_342; w_7_343<=Wgt_7_343; w_7_344<=Wgt_7_344; w_7_345<=Wgt_7_345; w_7_346<=Wgt_7_346; w_7_347<=Wgt_7_347; w_7_348<=Wgt_7_348; w_7_349<=Wgt_7_349; w_7_350<=Wgt_7_350; w_7_351<=Wgt_7_351; w_7_352<=Wgt_7_352; w_7_353<=Wgt_7_353; w_7_354<=Wgt_7_354; w_7_355<=Wgt_7_355; w_7_356<=Wgt_7_356; w_7_357<=Wgt_7_357; w_7_358<=Wgt_7_358; w_7_359<=Wgt_7_359; w_7_360<=Wgt_7_360; w_7_361<=Wgt_7_361; w_7_362<=Wgt_7_362; w_7_363<=Wgt_7_363; w_7_364<=Wgt_7_364; w_7_365<=Wgt_7_365; w_7_366<=Wgt_7_366; w_7_367<=Wgt_7_367; w_7_368<=Wgt_7_368; w_7_369<=Wgt_7_369; w_7_370<=Wgt_7_370; w_7_371<=Wgt_7_371; w_7_372<=Wgt_7_372; w_7_373<=Wgt_7_373; w_7_374<=Wgt_7_374; w_7_375<=Wgt_7_375; w_7_376<=Wgt_7_376; w_7_377<=Wgt_7_377; w_7_378<=Wgt_7_378; w_7_379<=Wgt_7_379; w_7_380<=Wgt_7_380; w_7_381<=Wgt_7_381; w_7_382<=Wgt_7_382; w_7_383<=Wgt_7_383; w_7_384<=Wgt_7_384; w_7_385<=Wgt_7_385; w_7_386<=Wgt_7_386; w_7_387<=Wgt_7_387; w_7_388<=Wgt_7_388; w_7_389<=Wgt_7_389; w_7_390<=Wgt_7_390; w_7_391<=Wgt_7_391; w_7_392<=Wgt_7_392; w_7_393<=Wgt_7_393; w_7_394<=Wgt_7_394; w_7_395<=Wgt_7_395; w_7_396<=Wgt_7_396; w_7_397<=Wgt_7_397; w_7_398<=Wgt_7_398; w_7_399<=Wgt_7_399; w_7_400<=Wgt_7_400; w_7_401<=Wgt_7_401; w_7_402<=Wgt_7_402; w_7_403<=Wgt_7_403; w_7_404<=Wgt_7_404; w_7_405<=Wgt_7_405; w_7_406<=Wgt_7_406; w_7_407<=Wgt_7_407; w_7_408<=Wgt_7_408; w_7_409<=Wgt_7_409; w_7_410<=Wgt_7_410; w_7_411<=Wgt_7_411; w_7_412<=Wgt_7_412; w_7_413<=Wgt_7_413; w_7_414<=Wgt_7_414; w_7_415<=Wgt_7_415; w_7_416<=Wgt_7_416; w_7_417<=Wgt_7_417; w_7_418<=Wgt_7_418; w_7_419<=Wgt_7_419; w_7_420<=Wgt_7_420; w_7_421<=Wgt_7_421; w_7_422<=Wgt_7_422; w_7_423<=Wgt_7_423; w_7_424<=Wgt_7_424; w_7_425<=Wgt_7_425; w_7_426<=Wgt_7_426; w_7_427<=Wgt_7_427; w_7_428<=Wgt_7_428; w_7_429<=Wgt_7_429; w_7_430<=Wgt_7_430; w_7_431<=Wgt_7_431; w_7_432<=Wgt_7_432; w_7_433<=Wgt_7_433; w_7_434<=Wgt_7_434; w_7_435<=Wgt_7_435; w_7_436<=Wgt_7_436; w_7_437<=Wgt_7_437; w_7_438<=Wgt_7_438; w_7_439<=Wgt_7_439; w_7_440<=Wgt_7_440; w_7_441<=Wgt_7_441; w_7_442<=Wgt_7_442; w_7_443<=Wgt_7_443; w_7_444<=Wgt_7_444; w_7_445<=Wgt_7_445; w_7_446<=Wgt_7_446; w_7_447<=Wgt_7_447; w_7_448<=Wgt_7_448; w_7_449<=Wgt_7_449; w_7_450<=Wgt_7_450; w_7_451<=Wgt_7_451; w_7_452<=Wgt_7_452; w_7_453<=Wgt_7_453; w_7_454<=Wgt_7_454; w_7_455<=Wgt_7_455; w_7_456<=Wgt_7_456; w_7_457<=Wgt_7_457; w_7_458<=Wgt_7_458; w_7_459<=Wgt_7_459; w_7_460<=Wgt_7_460; w_7_461<=Wgt_7_461; w_7_462<=Wgt_7_462; w_7_463<=Wgt_7_463; w_7_464<=Wgt_7_464; w_7_465<=Wgt_7_465; w_7_466<=Wgt_7_466; w_7_467<=Wgt_7_467; w_7_468<=Wgt_7_468; w_7_469<=Wgt_7_469; w_7_470<=Wgt_7_470; w_7_471<=Wgt_7_471; w_7_472<=Wgt_7_472; w_7_473<=Wgt_7_473; w_7_474<=Wgt_7_474; w_7_475<=Wgt_7_475; w_7_476<=Wgt_7_476; w_7_477<=Wgt_7_477; w_7_478<=Wgt_7_478; w_7_479<=Wgt_7_479; w_7_480<=Wgt_7_480; w_7_481<=Wgt_7_481; w_7_482<=Wgt_7_482; w_7_483<=Wgt_7_483; w_7_484<=Wgt_7_484; w_7_485<=Wgt_7_485; w_7_486<=Wgt_7_486; w_7_487<=Wgt_7_487; w_7_488<=Wgt_7_488; w_7_489<=Wgt_7_489; w_7_490<=Wgt_7_490; w_7_491<=Wgt_7_491; w_7_492<=Wgt_7_492; w_7_493<=Wgt_7_493; w_7_494<=Wgt_7_494; w_7_495<=Wgt_7_495; w_7_496<=Wgt_7_496; w_7_497<=Wgt_7_497; w_7_498<=Wgt_7_498; w_7_499<=Wgt_7_499; w_7_500<=Wgt_7_500; w_7_501<=Wgt_7_501; w_7_502<=Wgt_7_502; w_7_503<=Wgt_7_503; w_7_504<=Wgt_7_504; w_7_505<=Wgt_7_505; w_7_506<=Wgt_7_506; w_7_507<=Wgt_7_507; w_7_508<=Wgt_7_508; w_7_509<=Wgt_7_509; w_7_510<=Wgt_7_510; w_7_511<=Wgt_7_511; w_7_512<=Wgt_7_512; w_7_513<=Wgt_7_513; w_7_514<=Wgt_7_514; w_7_515<=Wgt_7_515; w_7_516<=Wgt_7_516; w_7_517<=Wgt_7_517; w_7_518<=Wgt_7_518; w_7_519<=Wgt_7_519; w_7_520<=Wgt_7_520; w_7_521<=Wgt_7_521; w_7_522<=Wgt_7_522; w_7_523<=Wgt_7_523; w_7_524<=Wgt_7_524; w_7_525<=Wgt_7_525; w_7_526<=Wgt_7_526; w_7_527<=Wgt_7_527; w_7_528<=Wgt_7_528; w_7_529<=Wgt_7_529; w_7_530<=Wgt_7_530; w_7_531<=Wgt_7_531; w_7_532<=Wgt_7_532; w_7_533<=Wgt_7_533; w_7_534<=Wgt_7_534; w_7_535<=Wgt_7_535; w_7_536<=Wgt_7_536; w_7_537<=Wgt_7_537; w_7_538<=Wgt_7_538; w_7_539<=Wgt_7_539; w_7_540<=Wgt_7_540; w_7_541<=Wgt_7_541; w_7_542<=Wgt_7_542; w_7_543<=Wgt_7_543; w_7_544<=Wgt_7_544; w_7_545<=Wgt_7_545; w_7_546<=Wgt_7_546; w_7_547<=Wgt_7_547; w_7_548<=Wgt_7_548; w_7_549<=Wgt_7_549; w_7_550<=Wgt_7_550; w_7_551<=Wgt_7_551; w_7_552<=Wgt_7_552; w_7_553<=Wgt_7_553; w_7_554<=Wgt_7_554; w_7_555<=Wgt_7_555; w_7_556<=Wgt_7_556; w_7_557<=Wgt_7_557; w_7_558<=Wgt_7_558; w_7_559<=Wgt_7_559; w_7_560<=Wgt_7_560; w_7_561<=Wgt_7_561; w_7_562<=Wgt_7_562; w_7_563<=Wgt_7_563; w_7_564<=Wgt_7_564; w_7_565<=Wgt_7_565; w_7_566<=Wgt_7_566; w_7_567<=Wgt_7_567; w_7_568<=Wgt_7_568; w_7_569<=Wgt_7_569; w_7_570<=Wgt_7_570; w_7_571<=Wgt_7_571; w_7_572<=Wgt_7_572; w_7_573<=Wgt_7_573; w_7_574<=Wgt_7_574; w_7_575<=Wgt_7_575; w_7_576<=Wgt_7_576; w_7_577<=Wgt_7_577; w_7_578<=Wgt_7_578; w_7_579<=Wgt_7_579; w_7_580<=Wgt_7_580; w_7_581<=Wgt_7_581; w_7_582<=Wgt_7_582; w_7_583<=Wgt_7_583; w_7_584<=Wgt_7_584; w_7_585<=Wgt_7_585; w_7_586<=Wgt_7_586; w_7_587<=Wgt_7_587; w_7_588<=Wgt_7_588; w_7_589<=Wgt_7_589; w_7_590<=Wgt_7_590; w_7_591<=Wgt_7_591; w_7_592<=Wgt_7_592; w_7_593<=Wgt_7_593; w_7_594<=Wgt_7_594; w_7_595<=Wgt_7_595; w_7_596<=Wgt_7_596; w_7_597<=Wgt_7_597; w_7_598<=Wgt_7_598; w_7_599<=Wgt_7_599; w_7_600<=Wgt_7_600; w_7_601<=Wgt_7_601; w_7_602<=Wgt_7_602; w_7_603<=Wgt_7_603; w_7_604<=Wgt_7_604; w_7_605<=Wgt_7_605; w_7_606<=Wgt_7_606; w_7_607<=Wgt_7_607; w_7_608<=Wgt_7_608; w_7_609<=Wgt_7_609; w_7_610<=Wgt_7_610; w_7_611<=Wgt_7_611; w_7_612<=Wgt_7_612; w_7_613<=Wgt_7_613; w_7_614<=Wgt_7_614; w_7_615<=Wgt_7_615; w_7_616<=Wgt_7_616; w_7_617<=Wgt_7_617; w_7_618<=Wgt_7_618; w_7_619<=Wgt_7_619; w_7_620<=Wgt_7_620; w_7_621<=Wgt_7_621; w_7_622<=Wgt_7_622; w_7_623<=Wgt_7_623; w_7_624<=Wgt_7_624; w_7_625<=Wgt_7_625; w_7_626<=Wgt_7_626; w_7_627<=Wgt_7_627; w_7_628<=Wgt_7_628; w_7_629<=Wgt_7_629; w_7_630<=Wgt_7_630; w_7_631<=Wgt_7_631; w_7_632<=Wgt_7_632; w_7_633<=Wgt_7_633; w_7_634<=Wgt_7_634; w_7_635<=Wgt_7_635; w_7_636<=Wgt_7_636; w_7_637<=Wgt_7_637; w_7_638<=Wgt_7_638; w_7_639<=Wgt_7_639; w_7_640<=Wgt_7_640; w_7_641<=Wgt_7_641; w_7_642<=Wgt_7_642; w_7_643<=Wgt_7_643; w_7_644<=Wgt_7_644; w_7_645<=Wgt_7_645; w_7_646<=Wgt_7_646; w_7_647<=Wgt_7_647; w_7_648<=Wgt_7_648; w_7_649<=Wgt_7_649; w_7_650<=Wgt_7_650; w_7_651<=Wgt_7_651; w_7_652<=Wgt_7_652; w_7_653<=Wgt_7_653; w_7_654<=Wgt_7_654; w_7_655<=Wgt_7_655; w_7_656<=Wgt_7_656; w_7_657<=Wgt_7_657; w_7_658<=Wgt_7_658; w_7_659<=Wgt_7_659; w_7_660<=Wgt_7_660; w_7_661<=Wgt_7_661; w_7_662<=Wgt_7_662; w_7_663<=Wgt_7_663; w_7_664<=Wgt_7_664; w_7_665<=Wgt_7_665; w_7_666<=Wgt_7_666; w_7_667<=Wgt_7_667; w_7_668<=Wgt_7_668; w_7_669<=Wgt_7_669; w_7_670<=Wgt_7_670; w_7_671<=Wgt_7_671; w_7_672<=Wgt_7_672; w_7_673<=Wgt_7_673; w_7_674<=Wgt_7_674; w_7_675<=Wgt_7_675; w_7_676<=Wgt_7_676; w_7_677<=Wgt_7_677; w_7_678<=Wgt_7_678; w_7_679<=Wgt_7_679; w_7_680<=Wgt_7_680; w_7_681<=Wgt_7_681; w_7_682<=Wgt_7_682; w_7_683<=Wgt_7_683; w_7_684<=Wgt_7_684; w_7_685<=Wgt_7_685; w_7_686<=Wgt_7_686; w_7_687<=Wgt_7_687; w_7_688<=Wgt_7_688; w_7_689<=Wgt_7_689; w_7_690<=Wgt_7_690; w_7_691<=Wgt_7_691; w_7_692<=Wgt_7_692; w_7_693<=Wgt_7_693; w_7_694<=Wgt_7_694; w_7_695<=Wgt_7_695; w_7_696<=Wgt_7_696; w_7_697<=Wgt_7_697; w_7_698<=Wgt_7_698; w_7_699<=Wgt_7_699; w_7_700<=Wgt_7_700; w_7_701<=Wgt_7_701; w_7_702<=Wgt_7_702; w_7_703<=Wgt_7_703; w_7_704<=Wgt_7_704; w_7_705<=Wgt_7_705; w_7_706<=Wgt_7_706; w_7_707<=Wgt_7_707; w_7_708<=Wgt_7_708; w_7_709<=Wgt_7_709; w_7_710<=Wgt_7_710; w_7_711<=Wgt_7_711; w_7_712<=Wgt_7_712; w_7_713<=Wgt_7_713; w_7_714<=Wgt_7_714; w_7_715<=Wgt_7_715; w_7_716<=Wgt_7_716; w_7_717<=Wgt_7_717; w_7_718<=Wgt_7_718; w_7_719<=Wgt_7_719; w_7_720<=Wgt_7_720; w_7_721<=Wgt_7_721; w_7_722<=Wgt_7_722; w_7_723<=Wgt_7_723; w_7_724<=Wgt_7_724; w_7_725<=Wgt_7_725; w_7_726<=Wgt_7_726; w_7_727<=Wgt_7_727; w_7_728<=Wgt_7_728; w_7_729<=Wgt_7_729; w_7_730<=Wgt_7_730; w_7_731<=Wgt_7_731; w_7_732<=Wgt_7_732; w_7_733<=Wgt_7_733; w_7_734<=Wgt_7_734; w_7_735<=Wgt_7_735; w_7_736<=Wgt_7_736; w_7_737<=Wgt_7_737; w_7_738<=Wgt_7_738; w_7_739<=Wgt_7_739; w_7_740<=Wgt_7_740; w_7_741<=Wgt_7_741; w_7_742<=Wgt_7_742; w_7_743<=Wgt_7_743; w_7_744<=Wgt_7_744; w_7_745<=Wgt_7_745; w_7_746<=Wgt_7_746; w_7_747<=Wgt_7_747; w_7_748<=Wgt_7_748; w_7_749<=Wgt_7_749; w_7_750<=Wgt_7_750; w_7_751<=Wgt_7_751; w_7_752<=Wgt_7_752; w_7_753<=Wgt_7_753; w_7_754<=Wgt_7_754; w_7_755<=Wgt_7_755; w_7_756<=Wgt_7_756; w_7_757<=Wgt_7_757; w_7_758<=Wgt_7_758; w_7_759<=Wgt_7_759; w_7_760<=Wgt_7_760; w_7_761<=Wgt_7_761; w_7_762<=Wgt_7_762; w_7_763<=Wgt_7_763; w_7_764<=Wgt_7_764; w_7_765<=Wgt_7_765; w_7_766<=Wgt_7_766; w_7_767<=Wgt_7_767; w_7_768<=Wgt_7_768; w_7_769<=Wgt_7_769; w_7_770<=Wgt_7_770; w_7_771<=Wgt_7_771; w_7_772<=Wgt_7_772; w_7_773<=Wgt_7_773; w_7_774<=Wgt_7_774; w_7_775<=Wgt_7_775; w_7_776<=Wgt_7_776; w_7_777<=Wgt_7_777; w_7_778<=Wgt_7_778; w_7_779<=Wgt_7_779; w_7_780<=Wgt_7_780; w_7_781<=Wgt_7_781; w_7_782<=Wgt_7_782; w_7_783<=Wgt_7_783; w_7_784<=Wgt_7_784; 
					w_8_0<=Wgt_8_0; w_8_1<=Wgt_8_1; w_8_2<=Wgt_8_2; w_8_3<=Wgt_8_3; w_8_4<=Wgt_8_4; w_8_5<=Wgt_8_5; w_8_6<=Wgt_8_6; w_8_7<=Wgt_8_7; w_8_8<=Wgt_8_8; w_8_9<=Wgt_8_9; w_8_10<=Wgt_8_10; w_8_11<=Wgt_8_11; w_8_12<=Wgt_8_12; w_8_13<=Wgt_8_13; w_8_14<=Wgt_8_14; w_8_15<=Wgt_8_15; w_8_16<=Wgt_8_16; w_8_17<=Wgt_8_17; w_8_18<=Wgt_8_18; w_8_19<=Wgt_8_19; w_8_20<=Wgt_8_20; w_8_21<=Wgt_8_21; w_8_22<=Wgt_8_22; w_8_23<=Wgt_8_23; w_8_24<=Wgt_8_24; w_8_25<=Wgt_8_25; w_8_26<=Wgt_8_26; w_8_27<=Wgt_8_27; w_8_28<=Wgt_8_28; w_8_29<=Wgt_8_29; w_8_30<=Wgt_8_30; w_8_31<=Wgt_8_31; w_8_32<=Wgt_8_32; w_8_33<=Wgt_8_33; w_8_34<=Wgt_8_34; w_8_35<=Wgt_8_35; w_8_36<=Wgt_8_36; w_8_37<=Wgt_8_37; w_8_38<=Wgt_8_38; w_8_39<=Wgt_8_39; w_8_40<=Wgt_8_40; w_8_41<=Wgt_8_41; w_8_42<=Wgt_8_42; w_8_43<=Wgt_8_43; w_8_44<=Wgt_8_44; w_8_45<=Wgt_8_45; w_8_46<=Wgt_8_46; w_8_47<=Wgt_8_47; w_8_48<=Wgt_8_48; w_8_49<=Wgt_8_49; w_8_50<=Wgt_8_50; w_8_51<=Wgt_8_51; w_8_52<=Wgt_8_52; w_8_53<=Wgt_8_53; w_8_54<=Wgt_8_54; w_8_55<=Wgt_8_55; w_8_56<=Wgt_8_56; w_8_57<=Wgt_8_57; w_8_58<=Wgt_8_58; w_8_59<=Wgt_8_59; w_8_60<=Wgt_8_60; w_8_61<=Wgt_8_61; w_8_62<=Wgt_8_62; w_8_63<=Wgt_8_63; w_8_64<=Wgt_8_64; w_8_65<=Wgt_8_65; w_8_66<=Wgt_8_66; w_8_67<=Wgt_8_67; w_8_68<=Wgt_8_68; w_8_69<=Wgt_8_69; w_8_70<=Wgt_8_70; w_8_71<=Wgt_8_71; w_8_72<=Wgt_8_72; w_8_73<=Wgt_8_73; w_8_74<=Wgt_8_74; w_8_75<=Wgt_8_75; w_8_76<=Wgt_8_76; w_8_77<=Wgt_8_77; w_8_78<=Wgt_8_78; w_8_79<=Wgt_8_79; w_8_80<=Wgt_8_80; w_8_81<=Wgt_8_81; w_8_82<=Wgt_8_82; w_8_83<=Wgt_8_83; w_8_84<=Wgt_8_84; w_8_85<=Wgt_8_85; w_8_86<=Wgt_8_86; w_8_87<=Wgt_8_87; w_8_88<=Wgt_8_88; w_8_89<=Wgt_8_89; w_8_90<=Wgt_8_90; w_8_91<=Wgt_8_91; w_8_92<=Wgt_8_92; w_8_93<=Wgt_8_93; w_8_94<=Wgt_8_94; w_8_95<=Wgt_8_95; w_8_96<=Wgt_8_96; w_8_97<=Wgt_8_97; w_8_98<=Wgt_8_98; w_8_99<=Wgt_8_99; w_8_100<=Wgt_8_100; w_8_101<=Wgt_8_101; w_8_102<=Wgt_8_102; w_8_103<=Wgt_8_103; w_8_104<=Wgt_8_104; w_8_105<=Wgt_8_105; w_8_106<=Wgt_8_106; w_8_107<=Wgt_8_107; w_8_108<=Wgt_8_108; w_8_109<=Wgt_8_109; w_8_110<=Wgt_8_110; w_8_111<=Wgt_8_111; w_8_112<=Wgt_8_112; w_8_113<=Wgt_8_113; w_8_114<=Wgt_8_114; w_8_115<=Wgt_8_115; w_8_116<=Wgt_8_116; w_8_117<=Wgt_8_117; w_8_118<=Wgt_8_118; w_8_119<=Wgt_8_119; w_8_120<=Wgt_8_120; w_8_121<=Wgt_8_121; w_8_122<=Wgt_8_122; w_8_123<=Wgt_8_123; w_8_124<=Wgt_8_124; w_8_125<=Wgt_8_125; w_8_126<=Wgt_8_126; w_8_127<=Wgt_8_127; w_8_128<=Wgt_8_128; w_8_129<=Wgt_8_129; w_8_130<=Wgt_8_130; w_8_131<=Wgt_8_131; w_8_132<=Wgt_8_132; w_8_133<=Wgt_8_133; w_8_134<=Wgt_8_134; w_8_135<=Wgt_8_135; w_8_136<=Wgt_8_136; w_8_137<=Wgt_8_137; w_8_138<=Wgt_8_138; w_8_139<=Wgt_8_139; w_8_140<=Wgt_8_140; w_8_141<=Wgt_8_141; w_8_142<=Wgt_8_142; w_8_143<=Wgt_8_143; w_8_144<=Wgt_8_144; w_8_145<=Wgt_8_145; w_8_146<=Wgt_8_146; w_8_147<=Wgt_8_147; w_8_148<=Wgt_8_148; w_8_149<=Wgt_8_149; w_8_150<=Wgt_8_150; w_8_151<=Wgt_8_151; w_8_152<=Wgt_8_152; w_8_153<=Wgt_8_153; w_8_154<=Wgt_8_154; w_8_155<=Wgt_8_155; w_8_156<=Wgt_8_156; w_8_157<=Wgt_8_157; w_8_158<=Wgt_8_158; w_8_159<=Wgt_8_159; w_8_160<=Wgt_8_160; w_8_161<=Wgt_8_161; w_8_162<=Wgt_8_162; w_8_163<=Wgt_8_163; w_8_164<=Wgt_8_164; w_8_165<=Wgt_8_165; w_8_166<=Wgt_8_166; w_8_167<=Wgt_8_167; w_8_168<=Wgt_8_168; w_8_169<=Wgt_8_169; w_8_170<=Wgt_8_170; w_8_171<=Wgt_8_171; w_8_172<=Wgt_8_172; w_8_173<=Wgt_8_173; w_8_174<=Wgt_8_174; w_8_175<=Wgt_8_175; w_8_176<=Wgt_8_176; w_8_177<=Wgt_8_177; w_8_178<=Wgt_8_178; w_8_179<=Wgt_8_179; w_8_180<=Wgt_8_180; w_8_181<=Wgt_8_181; w_8_182<=Wgt_8_182; w_8_183<=Wgt_8_183; w_8_184<=Wgt_8_184; w_8_185<=Wgt_8_185; w_8_186<=Wgt_8_186; w_8_187<=Wgt_8_187; w_8_188<=Wgt_8_188; w_8_189<=Wgt_8_189; w_8_190<=Wgt_8_190; w_8_191<=Wgt_8_191; w_8_192<=Wgt_8_192; w_8_193<=Wgt_8_193; w_8_194<=Wgt_8_194; w_8_195<=Wgt_8_195; w_8_196<=Wgt_8_196; w_8_197<=Wgt_8_197; w_8_198<=Wgt_8_198; w_8_199<=Wgt_8_199; w_8_200<=Wgt_8_200; w_8_201<=Wgt_8_201; w_8_202<=Wgt_8_202; w_8_203<=Wgt_8_203; w_8_204<=Wgt_8_204; w_8_205<=Wgt_8_205; w_8_206<=Wgt_8_206; w_8_207<=Wgt_8_207; w_8_208<=Wgt_8_208; w_8_209<=Wgt_8_209; w_8_210<=Wgt_8_210; w_8_211<=Wgt_8_211; w_8_212<=Wgt_8_212; w_8_213<=Wgt_8_213; w_8_214<=Wgt_8_214; w_8_215<=Wgt_8_215; w_8_216<=Wgt_8_216; w_8_217<=Wgt_8_217; w_8_218<=Wgt_8_218; w_8_219<=Wgt_8_219; w_8_220<=Wgt_8_220; w_8_221<=Wgt_8_221; w_8_222<=Wgt_8_222; w_8_223<=Wgt_8_223; w_8_224<=Wgt_8_224; w_8_225<=Wgt_8_225; w_8_226<=Wgt_8_226; w_8_227<=Wgt_8_227; w_8_228<=Wgt_8_228; w_8_229<=Wgt_8_229; w_8_230<=Wgt_8_230; w_8_231<=Wgt_8_231; w_8_232<=Wgt_8_232; w_8_233<=Wgt_8_233; w_8_234<=Wgt_8_234; w_8_235<=Wgt_8_235; w_8_236<=Wgt_8_236; w_8_237<=Wgt_8_237; w_8_238<=Wgt_8_238; w_8_239<=Wgt_8_239; w_8_240<=Wgt_8_240; w_8_241<=Wgt_8_241; w_8_242<=Wgt_8_242; w_8_243<=Wgt_8_243; w_8_244<=Wgt_8_244; w_8_245<=Wgt_8_245; w_8_246<=Wgt_8_246; w_8_247<=Wgt_8_247; w_8_248<=Wgt_8_248; w_8_249<=Wgt_8_249; w_8_250<=Wgt_8_250; w_8_251<=Wgt_8_251; w_8_252<=Wgt_8_252; w_8_253<=Wgt_8_253; w_8_254<=Wgt_8_254; w_8_255<=Wgt_8_255; w_8_256<=Wgt_8_256; w_8_257<=Wgt_8_257; w_8_258<=Wgt_8_258; w_8_259<=Wgt_8_259; w_8_260<=Wgt_8_260; w_8_261<=Wgt_8_261; w_8_262<=Wgt_8_262; w_8_263<=Wgt_8_263; w_8_264<=Wgt_8_264; w_8_265<=Wgt_8_265; w_8_266<=Wgt_8_266; w_8_267<=Wgt_8_267; w_8_268<=Wgt_8_268; w_8_269<=Wgt_8_269; w_8_270<=Wgt_8_270; w_8_271<=Wgt_8_271; w_8_272<=Wgt_8_272; w_8_273<=Wgt_8_273; w_8_274<=Wgt_8_274; w_8_275<=Wgt_8_275; w_8_276<=Wgt_8_276; w_8_277<=Wgt_8_277; w_8_278<=Wgt_8_278; w_8_279<=Wgt_8_279; w_8_280<=Wgt_8_280; w_8_281<=Wgt_8_281; w_8_282<=Wgt_8_282; w_8_283<=Wgt_8_283; w_8_284<=Wgt_8_284; w_8_285<=Wgt_8_285; w_8_286<=Wgt_8_286; w_8_287<=Wgt_8_287; w_8_288<=Wgt_8_288; w_8_289<=Wgt_8_289; w_8_290<=Wgt_8_290; w_8_291<=Wgt_8_291; w_8_292<=Wgt_8_292; w_8_293<=Wgt_8_293; w_8_294<=Wgt_8_294; w_8_295<=Wgt_8_295; w_8_296<=Wgt_8_296; w_8_297<=Wgt_8_297; w_8_298<=Wgt_8_298; w_8_299<=Wgt_8_299; w_8_300<=Wgt_8_300; w_8_301<=Wgt_8_301; w_8_302<=Wgt_8_302; w_8_303<=Wgt_8_303; w_8_304<=Wgt_8_304; w_8_305<=Wgt_8_305; w_8_306<=Wgt_8_306; w_8_307<=Wgt_8_307; w_8_308<=Wgt_8_308; w_8_309<=Wgt_8_309; w_8_310<=Wgt_8_310; w_8_311<=Wgt_8_311; w_8_312<=Wgt_8_312; w_8_313<=Wgt_8_313; w_8_314<=Wgt_8_314; w_8_315<=Wgt_8_315; w_8_316<=Wgt_8_316; w_8_317<=Wgt_8_317; w_8_318<=Wgt_8_318; w_8_319<=Wgt_8_319; w_8_320<=Wgt_8_320; w_8_321<=Wgt_8_321; w_8_322<=Wgt_8_322; w_8_323<=Wgt_8_323; w_8_324<=Wgt_8_324; w_8_325<=Wgt_8_325; w_8_326<=Wgt_8_326; w_8_327<=Wgt_8_327; w_8_328<=Wgt_8_328; w_8_329<=Wgt_8_329; w_8_330<=Wgt_8_330; w_8_331<=Wgt_8_331; w_8_332<=Wgt_8_332; w_8_333<=Wgt_8_333; w_8_334<=Wgt_8_334; w_8_335<=Wgt_8_335; w_8_336<=Wgt_8_336; w_8_337<=Wgt_8_337; w_8_338<=Wgt_8_338; w_8_339<=Wgt_8_339; w_8_340<=Wgt_8_340; w_8_341<=Wgt_8_341; w_8_342<=Wgt_8_342; w_8_343<=Wgt_8_343; w_8_344<=Wgt_8_344; w_8_345<=Wgt_8_345; w_8_346<=Wgt_8_346; w_8_347<=Wgt_8_347; w_8_348<=Wgt_8_348; w_8_349<=Wgt_8_349; w_8_350<=Wgt_8_350; w_8_351<=Wgt_8_351; w_8_352<=Wgt_8_352; w_8_353<=Wgt_8_353; w_8_354<=Wgt_8_354; w_8_355<=Wgt_8_355; w_8_356<=Wgt_8_356; w_8_357<=Wgt_8_357; w_8_358<=Wgt_8_358; w_8_359<=Wgt_8_359; w_8_360<=Wgt_8_360; w_8_361<=Wgt_8_361; w_8_362<=Wgt_8_362; w_8_363<=Wgt_8_363; w_8_364<=Wgt_8_364; w_8_365<=Wgt_8_365; w_8_366<=Wgt_8_366; w_8_367<=Wgt_8_367; w_8_368<=Wgt_8_368; w_8_369<=Wgt_8_369; w_8_370<=Wgt_8_370; w_8_371<=Wgt_8_371; w_8_372<=Wgt_8_372; w_8_373<=Wgt_8_373; w_8_374<=Wgt_8_374; w_8_375<=Wgt_8_375; w_8_376<=Wgt_8_376; w_8_377<=Wgt_8_377; w_8_378<=Wgt_8_378; w_8_379<=Wgt_8_379; w_8_380<=Wgt_8_380; w_8_381<=Wgt_8_381; w_8_382<=Wgt_8_382; w_8_383<=Wgt_8_383; w_8_384<=Wgt_8_384; w_8_385<=Wgt_8_385; w_8_386<=Wgt_8_386; w_8_387<=Wgt_8_387; w_8_388<=Wgt_8_388; w_8_389<=Wgt_8_389; w_8_390<=Wgt_8_390; w_8_391<=Wgt_8_391; w_8_392<=Wgt_8_392; w_8_393<=Wgt_8_393; w_8_394<=Wgt_8_394; w_8_395<=Wgt_8_395; w_8_396<=Wgt_8_396; w_8_397<=Wgt_8_397; w_8_398<=Wgt_8_398; w_8_399<=Wgt_8_399; w_8_400<=Wgt_8_400; w_8_401<=Wgt_8_401; w_8_402<=Wgt_8_402; w_8_403<=Wgt_8_403; w_8_404<=Wgt_8_404; w_8_405<=Wgt_8_405; w_8_406<=Wgt_8_406; w_8_407<=Wgt_8_407; w_8_408<=Wgt_8_408; w_8_409<=Wgt_8_409; w_8_410<=Wgt_8_410; w_8_411<=Wgt_8_411; w_8_412<=Wgt_8_412; w_8_413<=Wgt_8_413; w_8_414<=Wgt_8_414; w_8_415<=Wgt_8_415; w_8_416<=Wgt_8_416; w_8_417<=Wgt_8_417; w_8_418<=Wgt_8_418; w_8_419<=Wgt_8_419; w_8_420<=Wgt_8_420; w_8_421<=Wgt_8_421; w_8_422<=Wgt_8_422; w_8_423<=Wgt_8_423; w_8_424<=Wgt_8_424; w_8_425<=Wgt_8_425; w_8_426<=Wgt_8_426; w_8_427<=Wgt_8_427; w_8_428<=Wgt_8_428; w_8_429<=Wgt_8_429; w_8_430<=Wgt_8_430; w_8_431<=Wgt_8_431; w_8_432<=Wgt_8_432; w_8_433<=Wgt_8_433; w_8_434<=Wgt_8_434; w_8_435<=Wgt_8_435; w_8_436<=Wgt_8_436; w_8_437<=Wgt_8_437; w_8_438<=Wgt_8_438; w_8_439<=Wgt_8_439; w_8_440<=Wgt_8_440; w_8_441<=Wgt_8_441; w_8_442<=Wgt_8_442; w_8_443<=Wgt_8_443; w_8_444<=Wgt_8_444; w_8_445<=Wgt_8_445; w_8_446<=Wgt_8_446; w_8_447<=Wgt_8_447; w_8_448<=Wgt_8_448; w_8_449<=Wgt_8_449; w_8_450<=Wgt_8_450; w_8_451<=Wgt_8_451; w_8_452<=Wgt_8_452; w_8_453<=Wgt_8_453; w_8_454<=Wgt_8_454; w_8_455<=Wgt_8_455; w_8_456<=Wgt_8_456; w_8_457<=Wgt_8_457; w_8_458<=Wgt_8_458; w_8_459<=Wgt_8_459; w_8_460<=Wgt_8_460; w_8_461<=Wgt_8_461; w_8_462<=Wgt_8_462; w_8_463<=Wgt_8_463; w_8_464<=Wgt_8_464; w_8_465<=Wgt_8_465; w_8_466<=Wgt_8_466; w_8_467<=Wgt_8_467; w_8_468<=Wgt_8_468; w_8_469<=Wgt_8_469; w_8_470<=Wgt_8_470; w_8_471<=Wgt_8_471; w_8_472<=Wgt_8_472; w_8_473<=Wgt_8_473; w_8_474<=Wgt_8_474; w_8_475<=Wgt_8_475; w_8_476<=Wgt_8_476; w_8_477<=Wgt_8_477; w_8_478<=Wgt_8_478; w_8_479<=Wgt_8_479; w_8_480<=Wgt_8_480; w_8_481<=Wgt_8_481; w_8_482<=Wgt_8_482; w_8_483<=Wgt_8_483; w_8_484<=Wgt_8_484; w_8_485<=Wgt_8_485; w_8_486<=Wgt_8_486; w_8_487<=Wgt_8_487; w_8_488<=Wgt_8_488; w_8_489<=Wgt_8_489; w_8_490<=Wgt_8_490; w_8_491<=Wgt_8_491; w_8_492<=Wgt_8_492; w_8_493<=Wgt_8_493; w_8_494<=Wgt_8_494; w_8_495<=Wgt_8_495; w_8_496<=Wgt_8_496; w_8_497<=Wgt_8_497; w_8_498<=Wgt_8_498; w_8_499<=Wgt_8_499; w_8_500<=Wgt_8_500; w_8_501<=Wgt_8_501; w_8_502<=Wgt_8_502; w_8_503<=Wgt_8_503; w_8_504<=Wgt_8_504; w_8_505<=Wgt_8_505; w_8_506<=Wgt_8_506; w_8_507<=Wgt_8_507; w_8_508<=Wgt_8_508; w_8_509<=Wgt_8_509; w_8_510<=Wgt_8_510; w_8_511<=Wgt_8_511; w_8_512<=Wgt_8_512; w_8_513<=Wgt_8_513; w_8_514<=Wgt_8_514; w_8_515<=Wgt_8_515; w_8_516<=Wgt_8_516; w_8_517<=Wgt_8_517; w_8_518<=Wgt_8_518; w_8_519<=Wgt_8_519; w_8_520<=Wgt_8_520; w_8_521<=Wgt_8_521; w_8_522<=Wgt_8_522; w_8_523<=Wgt_8_523; w_8_524<=Wgt_8_524; w_8_525<=Wgt_8_525; w_8_526<=Wgt_8_526; w_8_527<=Wgt_8_527; w_8_528<=Wgt_8_528; w_8_529<=Wgt_8_529; w_8_530<=Wgt_8_530; w_8_531<=Wgt_8_531; w_8_532<=Wgt_8_532; w_8_533<=Wgt_8_533; w_8_534<=Wgt_8_534; w_8_535<=Wgt_8_535; w_8_536<=Wgt_8_536; w_8_537<=Wgt_8_537; w_8_538<=Wgt_8_538; w_8_539<=Wgt_8_539; w_8_540<=Wgt_8_540; w_8_541<=Wgt_8_541; w_8_542<=Wgt_8_542; w_8_543<=Wgt_8_543; w_8_544<=Wgt_8_544; w_8_545<=Wgt_8_545; w_8_546<=Wgt_8_546; w_8_547<=Wgt_8_547; w_8_548<=Wgt_8_548; w_8_549<=Wgt_8_549; w_8_550<=Wgt_8_550; w_8_551<=Wgt_8_551; w_8_552<=Wgt_8_552; w_8_553<=Wgt_8_553; w_8_554<=Wgt_8_554; w_8_555<=Wgt_8_555; w_8_556<=Wgt_8_556; w_8_557<=Wgt_8_557; w_8_558<=Wgt_8_558; w_8_559<=Wgt_8_559; w_8_560<=Wgt_8_560; w_8_561<=Wgt_8_561; w_8_562<=Wgt_8_562; w_8_563<=Wgt_8_563; w_8_564<=Wgt_8_564; w_8_565<=Wgt_8_565; w_8_566<=Wgt_8_566; w_8_567<=Wgt_8_567; w_8_568<=Wgt_8_568; w_8_569<=Wgt_8_569; w_8_570<=Wgt_8_570; w_8_571<=Wgt_8_571; w_8_572<=Wgt_8_572; w_8_573<=Wgt_8_573; w_8_574<=Wgt_8_574; w_8_575<=Wgt_8_575; w_8_576<=Wgt_8_576; w_8_577<=Wgt_8_577; w_8_578<=Wgt_8_578; w_8_579<=Wgt_8_579; w_8_580<=Wgt_8_580; w_8_581<=Wgt_8_581; w_8_582<=Wgt_8_582; w_8_583<=Wgt_8_583; w_8_584<=Wgt_8_584; w_8_585<=Wgt_8_585; w_8_586<=Wgt_8_586; w_8_587<=Wgt_8_587; w_8_588<=Wgt_8_588; w_8_589<=Wgt_8_589; w_8_590<=Wgt_8_590; w_8_591<=Wgt_8_591; w_8_592<=Wgt_8_592; w_8_593<=Wgt_8_593; w_8_594<=Wgt_8_594; w_8_595<=Wgt_8_595; w_8_596<=Wgt_8_596; w_8_597<=Wgt_8_597; w_8_598<=Wgt_8_598; w_8_599<=Wgt_8_599; w_8_600<=Wgt_8_600; w_8_601<=Wgt_8_601; w_8_602<=Wgt_8_602; w_8_603<=Wgt_8_603; w_8_604<=Wgt_8_604; w_8_605<=Wgt_8_605; w_8_606<=Wgt_8_606; w_8_607<=Wgt_8_607; w_8_608<=Wgt_8_608; w_8_609<=Wgt_8_609; w_8_610<=Wgt_8_610; w_8_611<=Wgt_8_611; w_8_612<=Wgt_8_612; w_8_613<=Wgt_8_613; w_8_614<=Wgt_8_614; w_8_615<=Wgt_8_615; w_8_616<=Wgt_8_616; w_8_617<=Wgt_8_617; w_8_618<=Wgt_8_618; w_8_619<=Wgt_8_619; w_8_620<=Wgt_8_620; w_8_621<=Wgt_8_621; w_8_622<=Wgt_8_622; w_8_623<=Wgt_8_623; w_8_624<=Wgt_8_624; w_8_625<=Wgt_8_625; w_8_626<=Wgt_8_626; w_8_627<=Wgt_8_627; w_8_628<=Wgt_8_628; w_8_629<=Wgt_8_629; w_8_630<=Wgt_8_630; w_8_631<=Wgt_8_631; w_8_632<=Wgt_8_632; w_8_633<=Wgt_8_633; w_8_634<=Wgt_8_634; w_8_635<=Wgt_8_635; w_8_636<=Wgt_8_636; w_8_637<=Wgt_8_637; w_8_638<=Wgt_8_638; w_8_639<=Wgt_8_639; w_8_640<=Wgt_8_640; w_8_641<=Wgt_8_641; w_8_642<=Wgt_8_642; w_8_643<=Wgt_8_643; w_8_644<=Wgt_8_644; w_8_645<=Wgt_8_645; w_8_646<=Wgt_8_646; w_8_647<=Wgt_8_647; w_8_648<=Wgt_8_648; w_8_649<=Wgt_8_649; w_8_650<=Wgt_8_650; w_8_651<=Wgt_8_651; w_8_652<=Wgt_8_652; w_8_653<=Wgt_8_653; w_8_654<=Wgt_8_654; w_8_655<=Wgt_8_655; w_8_656<=Wgt_8_656; w_8_657<=Wgt_8_657; w_8_658<=Wgt_8_658; w_8_659<=Wgt_8_659; w_8_660<=Wgt_8_660; w_8_661<=Wgt_8_661; w_8_662<=Wgt_8_662; w_8_663<=Wgt_8_663; w_8_664<=Wgt_8_664; w_8_665<=Wgt_8_665; w_8_666<=Wgt_8_666; w_8_667<=Wgt_8_667; w_8_668<=Wgt_8_668; w_8_669<=Wgt_8_669; w_8_670<=Wgt_8_670; w_8_671<=Wgt_8_671; w_8_672<=Wgt_8_672; w_8_673<=Wgt_8_673; w_8_674<=Wgt_8_674; w_8_675<=Wgt_8_675; w_8_676<=Wgt_8_676; w_8_677<=Wgt_8_677; w_8_678<=Wgt_8_678; w_8_679<=Wgt_8_679; w_8_680<=Wgt_8_680; w_8_681<=Wgt_8_681; w_8_682<=Wgt_8_682; w_8_683<=Wgt_8_683; w_8_684<=Wgt_8_684; w_8_685<=Wgt_8_685; w_8_686<=Wgt_8_686; w_8_687<=Wgt_8_687; w_8_688<=Wgt_8_688; w_8_689<=Wgt_8_689; w_8_690<=Wgt_8_690; w_8_691<=Wgt_8_691; w_8_692<=Wgt_8_692; w_8_693<=Wgt_8_693; w_8_694<=Wgt_8_694; w_8_695<=Wgt_8_695; w_8_696<=Wgt_8_696; w_8_697<=Wgt_8_697; w_8_698<=Wgt_8_698; w_8_699<=Wgt_8_699; w_8_700<=Wgt_8_700; w_8_701<=Wgt_8_701; w_8_702<=Wgt_8_702; w_8_703<=Wgt_8_703; w_8_704<=Wgt_8_704; w_8_705<=Wgt_8_705; w_8_706<=Wgt_8_706; w_8_707<=Wgt_8_707; w_8_708<=Wgt_8_708; w_8_709<=Wgt_8_709; w_8_710<=Wgt_8_710; w_8_711<=Wgt_8_711; w_8_712<=Wgt_8_712; w_8_713<=Wgt_8_713; w_8_714<=Wgt_8_714; w_8_715<=Wgt_8_715; w_8_716<=Wgt_8_716; w_8_717<=Wgt_8_717; w_8_718<=Wgt_8_718; w_8_719<=Wgt_8_719; w_8_720<=Wgt_8_720; w_8_721<=Wgt_8_721; w_8_722<=Wgt_8_722; w_8_723<=Wgt_8_723; w_8_724<=Wgt_8_724; w_8_725<=Wgt_8_725; w_8_726<=Wgt_8_726; w_8_727<=Wgt_8_727; w_8_728<=Wgt_8_728; w_8_729<=Wgt_8_729; w_8_730<=Wgt_8_730; w_8_731<=Wgt_8_731; w_8_732<=Wgt_8_732; w_8_733<=Wgt_8_733; w_8_734<=Wgt_8_734; w_8_735<=Wgt_8_735; w_8_736<=Wgt_8_736; w_8_737<=Wgt_8_737; w_8_738<=Wgt_8_738; w_8_739<=Wgt_8_739; w_8_740<=Wgt_8_740; w_8_741<=Wgt_8_741; w_8_742<=Wgt_8_742; w_8_743<=Wgt_8_743; w_8_744<=Wgt_8_744; w_8_745<=Wgt_8_745; w_8_746<=Wgt_8_746; w_8_747<=Wgt_8_747; w_8_748<=Wgt_8_748; w_8_749<=Wgt_8_749; w_8_750<=Wgt_8_750; w_8_751<=Wgt_8_751; w_8_752<=Wgt_8_752; w_8_753<=Wgt_8_753; w_8_754<=Wgt_8_754; w_8_755<=Wgt_8_755; w_8_756<=Wgt_8_756; w_8_757<=Wgt_8_757; w_8_758<=Wgt_8_758; w_8_759<=Wgt_8_759; w_8_760<=Wgt_8_760; w_8_761<=Wgt_8_761; w_8_762<=Wgt_8_762; w_8_763<=Wgt_8_763; w_8_764<=Wgt_8_764; w_8_765<=Wgt_8_765; w_8_766<=Wgt_8_766; w_8_767<=Wgt_8_767; w_8_768<=Wgt_8_768; w_8_769<=Wgt_8_769; w_8_770<=Wgt_8_770; w_8_771<=Wgt_8_771; w_8_772<=Wgt_8_772; w_8_773<=Wgt_8_773; w_8_774<=Wgt_8_774; w_8_775<=Wgt_8_775; w_8_776<=Wgt_8_776; w_8_777<=Wgt_8_777; w_8_778<=Wgt_8_778; w_8_779<=Wgt_8_779; w_8_780<=Wgt_8_780; w_8_781<=Wgt_8_781; w_8_782<=Wgt_8_782; w_8_783<=Wgt_8_783; w_8_784<=Wgt_8_784; 
					w_9_0<=Wgt_9_0; w_9_1<=Wgt_9_1; w_9_2<=Wgt_9_2; w_9_3<=Wgt_9_3; w_9_4<=Wgt_9_4; w_9_5<=Wgt_9_5; w_9_6<=Wgt_9_6; w_9_7<=Wgt_9_7; w_9_8<=Wgt_9_8; w_9_9<=Wgt_9_9; w_9_10<=Wgt_9_10; w_9_11<=Wgt_9_11; w_9_12<=Wgt_9_12; w_9_13<=Wgt_9_13; w_9_14<=Wgt_9_14; w_9_15<=Wgt_9_15; w_9_16<=Wgt_9_16; w_9_17<=Wgt_9_17; w_9_18<=Wgt_9_18; w_9_19<=Wgt_9_19; w_9_20<=Wgt_9_20; w_9_21<=Wgt_9_21; w_9_22<=Wgt_9_22; w_9_23<=Wgt_9_23; w_9_24<=Wgt_9_24; w_9_25<=Wgt_9_25; w_9_26<=Wgt_9_26; w_9_27<=Wgt_9_27; w_9_28<=Wgt_9_28; w_9_29<=Wgt_9_29; w_9_30<=Wgt_9_30; w_9_31<=Wgt_9_31; w_9_32<=Wgt_9_32; w_9_33<=Wgt_9_33; w_9_34<=Wgt_9_34; w_9_35<=Wgt_9_35; w_9_36<=Wgt_9_36; w_9_37<=Wgt_9_37; w_9_38<=Wgt_9_38; w_9_39<=Wgt_9_39; w_9_40<=Wgt_9_40; w_9_41<=Wgt_9_41; w_9_42<=Wgt_9_42; w_9_43<=Wgt_9_43; w_9_44<=Wgt_9_44; w_9_45<=Wgt_9_45; w_9_46<=Wgt_9_46; w_9_47<=Wgt_9_47; w_9_48<=Wgt_9_48; w_9_49<=Wgt_9_49; w_9_50<=Wgt_9_50; w_9_51<=Wgt_9_51; w_9_52<=Wgt_9_52; w_9_53<=Wgt_9_53; w_9_54<=Wgt_9_54; w_9_55<=Wgt_9_55; w_9_56<=Wgt_9_56; w_9_57<=Wgt_9_57; w_9_58<=Wgt_9_58; w_9_59<=Wgt_9_59; w_9_60<=Wgt_9_60; w_9_61<=Wgt_9_61; w_9_62<=Wgt_9_62; w_9_63<=Wgt_9_63; w_9_64<=Wgt_9_64; w_9_65<=Wgt_9_65; w_9_66<=Wgt_9_66; w_9_67<=Wgt_9_67; w_9_68<=Wgt_9_68; w_9_69<=Wgt_9_69; w_9_70<=Wgt_9_70; w_9_71<=Wgt_9_71; w_9_72<=Wgt_9_72; w_9_73<=Wgt_9_73; w_9_74<=Wgt_9_74; w_9_75<=Wgt_9_75; w_9_76<=Wgt_9_76; w_9_77<=Wgt_9_77; w_9_78<=Wgt_9_78; w_9_79<=Wgt_9_79; w_9_80<=Wgt_9_80; w_9_81<=Wgt_9_81; w_9_82<=Wgt_9_82; w_9_83<=Wgt_9_83; w_9_84<=Wgt_9_84; w_9_85<=Wgt_9_85; w_9_86<=Wgt_9_86; w_9_87<=Wgt_9_87; w_9_88<=Wgt_9_88; w_9_89<=Wgt_9_89; w_9_90<=Wgt_9_90; w_9_91<=Wgt_9_91; w_9_92<=Wgt_9_92; w_9_93<=Wgt_9_93; w_9_94<=Wgt_9_94; w_9_95<=Wgt_9_95; w_9_96<=Wgt_9_96; w_9_97<=Wgt_9_97; w_9_98<=Wgt_9_98; w_9_99<=Wgt_9_99; w_9_100<=Wgt_9_100; w_9_101<=Wgt_9_101; w_9_102<=Wgt_9_102; w_9_103<=Wgt_9_103; w_9_104<=Wgt_9_104; w_9_105<=Wgt_9_105; w_9_106<=Wgt_9_106; w_9_107<=Wgt_9_107; w_9_108<=Wgt_9_108; w_9_109<=Wgt_9_109; w_9_110<=Wgt_9_110; w_9_111<=Wgt_9_111; w_9_112<=Wgt_9_112; w_9_113<=Wgt_9_113; w_9_114<=Wgt_9_114; w_9_115<=Wgt_9_115; w_9_116<=Wgt_9_116; w_9_117<=Wgt_9_117; w_9_118<=Wgt_9_118; w_9_119<=Wgt_9_119; w_9_120<=Wgt_9_120; w_9_121<=Wgt_9_121; w_9_122<=Wgt_9_122; w_9_123<=Wgt_9_123; w_9_124<=Wgt_9_124; w_9_125<=Wgt_9_125; w_9_126<=Wgt_9_126; w_9_127<=Wgt_9_127; w_9_128<=Wgt_9_128; w_9_129<=Wgt_9_129; w_9_130<=Wgt_9_130; w_9_131<=Wgt_9_131; w_9_132<=Wgt_9_132; w_9_133<=Wgt_9_133; w_9_134<=Wgt_9_134; w_9_135<=Wgt_9_135; w_9_136<=Wgt_9_136; w_9_137<=Wgt_9_137; w_9_138<=Wgt_9_138; w_9_139<=Wgt_9_139; w_9_140<=Wgt_9_140; w_9_141<=Wgt_9_141; w_9_142<=Wgt_9_142; w_9_143<=Wgt_9_143; w_9_144<=Wgt_9_144; w_9_145<=Wgt_9_145; w_9_146<=Wgt_9_146; w_9_147<=Wgt_9_147; w_9_148<=Wgt_9_148; w_9_149<=Wgt_9_149; w_9_150<=Wgt_9_150; w_9_151<=Wgt_9_151; w_9_152<=Wgt_9_152; w_9_153<=Wgt_9_153; w_9_154<=Wgt_9_154; w_9_155<=Wgt_9_155; w_9_156<=Wgt_9_156; w_9_157<=Wgt_9_157; w_9_158<=Wgt_9_158; w_9_159<=Wgt_9_159; w_9_160<=Wgt_9_160; w_9_161<=Wgt_9_161; w_9_162<=Wgt_9_162; w_9_163<=Wgt_9_163; w_9_164<=Wgt_9_164; w_9_165<=Wgt_9_165; w_9_166<=Wgt_9_166; w_9_167<=Wgt_9_167; w_9_168<=Wgt_9_168; w_9_169<=Wgt_9_169; w_9_170<=Wgt_9_170; w_9_171<=Wgt_9_171; w_9_172<=Wgt_9_172; w_9_173<=Wgt_9_173; w_9_174<=Wgt_9_174; w_9_175<=Wgt_9_175; w_9_176<=Wgt_9_176; w_9_177<=Wgt_9_177; w_9_178<=Wgt_9_178; w_9_179<=Wgt_9_179; w_9_180<=Wgt_9_180; w_9_181<=Wgt_9_181; w_9_182<=Wgt_9_182; w_9_183<=Wgt_9_183; w_9_184<=Wgt_9_184; w_9_185<=Wgt_9_185; w_9_186<=Wgt_9_186; w_9_187<=Wgt_9_187; w_9_188<=Wgt_9_188; w_9_189<=Wgt_9_189; w_9_190<=Wgt_9_190; w_9_191<=Wgt_9_191; w_9_192<=Wgt_9_192; w_9_193<=Wgt_9_193; w_9_194<=Wgt_9_194; w_9_195<=Wgt_9_195; w_9_196<=Wgt_9_196; w_9_197<=Wgt_9_197; w_9_198<=Wgt_9_198; w_9_199<=Wgt_9_199; w_9_200<=Wgt_9_200; w_9_201<=Wgt_9_201; w_9_202<=Wgt_9_202; w_9_203<=Wgt_9_203; w_9_204<=Wgt_9_204; w_9_205<=Wgt_9_205; w_9_206<=Wgt_9_206; w_9_207<=Wgt_9_207; w_9_208<=Wgt_9_208; w_9_209<=Wgt_9_209; w_9_210<=Wgt_9_210; w_9_211<=Wgt_9_211; w_9_212<=Wgt_9_212; w_9_213<=Wgt_9_213; w_9_214<=Wgt_9_214; w_9_215<=Wgt_9_215; w_9_216<=Wgt_9_216; w_9_217<=Wgt_9_217; w_9_218<=Wgt_9_218; w_9_219<=Wgt_9_219; w_9_220<=Wgt_9_220; w_9_221<=Wgt_9_221; w_9_222<=Wgt_9_222; w_9_223<=Wgt_9_223; w_9_224<=Wgt_9_224; w_9_225<=Wgt_9_225; w_9_226<=Wgt_9_226; w_9_227<=Wgt_9_227; w_9_228<=Wgt_9_228; w_9_229<=Wgt_9_229; w_9_230<=Wgt_9_230; w_9_231<=Wgt_9_231; w_9_232<=Wgt_9_232; w_9_233<=Wgt_9_233; w_9_234<=Wgt_9_234; w_9_235<=Wgt_9_235; w_9_236<=Wgt_9_236; w_9_237<=Wgt_9_237; w_9_238<=Wgt_9_238; w_9_239<=Wgt_9_239; w_9_240<=Wgt_9_240; w_9_241<=Wgt_9_241; w_9_242<=Wgt_9_242; w_9_243<=Wgt_9_243; w_9_244<=Wgt_9_244; w_9_245<=Wgt_9_245; w_9_246<=Wgt_9_246; w_9_247<=Wgt_9_247; w_9_248<=Wgt_9_248; w_9_249<=Wgt_9_249; w_9_250<=Wgt_9_250; w_9_251<=Wgt_9_251; w_9_252<=Wgt_9_252; w_9_253<=Wgt_9_253; w_9_254<=Wgt_9_254; w_9_255<=Wgt_9_255; w_9_256<=Wgt_9_256; w_9_257<=Wgt_9_257; w_9_258<=Wgt_9_258; w_9_259<=Wgt_9_259; w_9_260<=Wgt_9_260; w_9_261<=Wgt_9_261; w_9_262<=Wgt_9_262; w_9_263<=Wgt_9_263; w_9_264<=Wgt_9_264; w_9_265<=Wgt_9_265; w_9_266<=Wgt_9_266; w_9_267<=Wgt_9_267; w_9_268<=Wgt_9_268; w_9_269<=Wgt_9_269; w_9_270<=Wgt_9_270; w_9_271<=Wgt_9_271; w_9_272<=Wgt_9_272; w_9_273<=Wgt_9_273; w_9_274<=Wgt_9_274; w_9_275<=Wgt_9_275; w_9_276<=Wgt_9_276; w_9_277<=Wgt_9_277; w_9_278<=Wgt_9_278; w_9_279<=Wgt_9_279; w_9_280<=Wgt_9_280; w_9_281<=Wgt_9_281; w_9_282<=Wgt_9_282; w_9_283<=Wgt_9_283; w_9_284<=Wgt_9_284; w_9_285<=Wgt_9_285; w_9_286<=Wgt_9_286; w_9_287<=Wgt_9_287; w_9_288<=Wgt_9_288; w_9_289<=Wgt_9_289; w_9_290<=Wgt_9_290; w_9_291<=Wgt_9_291; w_9_292<=Wgt_9_292; w_9_293<=Wgt_9_293; w_9_294<=Wgt_9_294; w_9_295<=Wgt_9_295; w_9_296<=Wgt_9_296; w_9_297<=Wgt_9_297; w_9_298<=Wgt_9_298; w_9_299<=Wgt_9_299; w_9_300<=Wgt_9_300; w_9_301<=Wgt_9_301; w_9_302<=Wgt_9_302; w_9_303<=Wgt_9_303; w_9_304<=Wgt_9_304; w_9_305<=Wgt_9_305; w_9_306<=Wgt_9_306; w_9_307<=Wgt_9_307; w_9_308<=Wgt_9_308; w_9_309<=Wgt_9_309; w_9_310<=Wgt_9_310; w_9_311<=Wgt_9_311; w_9_312<=Wgt_9_312; w_9_313<=Wgt_9_313; w_9_314<=Wgt_9_314; w_9_315<=Wgt_9_315; w_9_316<=Wgt_9_316; w_9_317<=Wgt_9_317; w_9_318<=Wgt_9_318; w_9_319<=Wgt_9_319; w_9_320<=Wgt_9_320; w_9_321<=Wgt_9_321; w_9_322<=Wgt_9_322; w_9_323<=Wgt_9_323; w_9_324<=Wgt_9_324; w_9_325<=Wgt_9_325; w_9_326<=Wgt_9_326; w_9_327<=Wgt_9_327; w_9_328<=Wgt_9_328; w_9_329<=Wgt_9_329; w_9_330<=Wgt_9_330; w_9_331<=Wgt_9_331; w_9_332<=Wgt_9_332; w_9_333<=Wgt_9_333; w_9_334<=Wgt_9_334; w_9_335<=Wgt_9_335; w_9_336<=Wgt_9_336; w_9_337<=Wgt_9_337; w_9_338<=Wgt_9_338; w_9_339<=Wgt_9_339; w_9_340<=Wgt_9_340; w_9_341<=Wgt_9_341; w_9_342<=Wgt_9_342; w_9_343<=Wgt_9_343; w_9_344<=Wgt_9_344; w_9_345<=Wgt_9_345; w_9_346<=Wgt_9_346; w_9_347<=Wgt_9_347; w_9_348<=Wgt_9_348; w_9_349<=Wgt_9_349; w_9_350<=Wgt_9_350; w_9_351<=Wgt_9_351; w_9_352<=Wgt_9_352; w_9_353<=Wgt_9_353; w_9_354<=Wgt_9_354; w_9_355<=Wgt_9_355; w_9_356<=Wgt_9_356; w_9_357<=Wgt_9_357; w_9_358<=Wgt_9_358; w_9_359<=Wgt_9_359; w_9_360<=Wgt_9_360; w_9_361<=Wgt_9_361; w_9_362<=Wgt_9_362; w_9_363<=Wgt_9_363; w_9_364<=Wgt_9_364; w_9_365<=Wgt_9_365; w_9_366<=Wgt_9_366; w_9_367<=Wgt_9_367; w_9_368<=Wgt_9_368; w_9_369<=Wgt_9_369; w_9_370<=Wgt_9_370; w_9_371<=Wgt_9_371; w_9_372<=Wgt_9_372; w_9_373<=Wgt_9_373; w_9_374<=Wgt_9_374; w_9_375<=Wgt_9_375; w_9_376<=Wgt_9_376; w_9_377<=Wgt_9_377; w_9_378<=Wgt_9_378; w_9_379<=Wgt_9_379; w_9_380<=Wgt_9_380; w_9_381<=Wgt_9_381; w_9_382<=Wgt_9_382; w_9_383<=Wgt_9_383; w_9_384<=Wgt_9_384; w_9_385<=Wgt_9_385; w_9_386<=Wgt_9_386; w_9_387<=Wgt_9_387; w_9_388<=Wgt_9_388; w_9_389<=Wgt_9_389; w_9_390<=Wgt_9_390; w_9_391<=Wgt_9_391; w_9_392<=Wgt_9_392; w_9_393<=Wgt_9_393; w_9_394<=Wgt_9_394; w_9_395<=Wgt_9_395; w_9_396<=Wgt_9_396; w_9_397<=Wgt_9_397; w_9_398<=Wgt_9_398; w_9_399<=Wgt_9_399; w_9_400<=Wgt_9_400; w_9_401<=Wgt_9_401; w_9_402<=Wgt_9_402; w_9_403<=Wgt_9_403; w_9_404<=Wgt_9_404; w_9_405<=Wgt_9_405; w_9_406<=Wgt_9_406; w_9_407<=Wgt_9_407; w_9_408<=Wgt_9_408; w_9_409<=Wgt_9_409; w_9_410<=Wgt_9_410; w_9_411<=Wgt_9_411; w_9_412<=Wgt_9_412; w_9_413<=Wgt_9_413; w_9_414<=Wgt_9_414; w_9_415<=Wgt_9_415; w_9_416<=Wgt_9_416; w_9_417<=Wgt_9_417; w_9_418<=Wgt_9_418; w_9_419<=Wgt_9_419; w_9_420<=Wgt_9_420; w_9_421<=Wgt_9_421; w_9_422<=Wgt_9_422; w_9_423<=Wgt_9_423; w_9_424<=Wgt_9_424; w_9_425<=Wgt_9_425; w_9_426<=Wgt_9_426; w_9_427<=Wgt_9_427; w_9_428<=Wgt_9_428; w_9_429<=Wgt_9_429; w_9_430<=Wgt_9_430; w_9_431<=Wgt_9_431; w_9_432<=Wgt_9_432; w_9_433<=Wgt_9_433; w_9_434<=Wgt_9_434; w_9_435<=Wgt_9_435; w_9_436<=Wgt_9_436; w_9_437<=Wgt_9_437; w_9_438<=Wgt_9_438; w_9_439<=Wgt_9_439; w_9_440<=Wgt_9_440; w_9_441<=Wgt_9_441; w_9_442<=Wgt_9_442; w_9_443<=Wgt_9_443; w_9_444<=Wgt_9_444; w_9_445<=Wgt_9_445; w_9_446<=Wgt_9_446; w_9_447<=Wgt_9_447; w_9_448<=Wgt_9_448; w_9_449<=Wgt_9_449; w_9_450<=Wgt_9_450; w_9_451<=Wgt_9_451; w_9_452<=Wgt_9_452; w_9_453<=Wgt_9_453; w_9_454<=Wgt_9_454; w_9_455<=Wgt_9_455; w_9_456<=Wgt_9_456; w_9_457<=Wgt_9_457; w_9_458<=Wgt_9_458; w_9_459<=Wgt_9_459; w_9_460<=Wgt_9_460; w_9_461<=Wgt_9_461; w_9_462<=Wgt_9_462; w_9_463<=Wgt_9_463; w_9_464<=Wgt_9_464; w_9_465<=Wgt_9_465; w_9_466<=Wgt_9_466; w_9_467<=Wgt_9_467; w_9_468<=Wgt_9_468; w_9_469<=Wgt_9_469; w_9_470<=Wgt_9_470; w_9_471<=Wgt_9_471; w_9_472<=Wgt_9_472; w_9_473<=Wgt_9_473; w_9_474<=Wgt_9_474; w_9_475<=Wgt_9_475; w_9_476<=Wgt_9_476; w_9_477<=Wgt_9_477; w_9_478<=Wgt_9_478; w_9_479<=Wgt_9_479; w_9_480<=Wgt_9_480; w_9_481<=Wgt_9_481; w_9_482<=Wgt_9_482; w_9_483<=Wgt_9_483; w_9_484<=Wgt_9_484; w_9_485<=Wgt_9_485; w_9_486<=Wgt_9_486; w_9_487<=Wgt_9_487; w_9_488<=Wgt_9_488; w_9_489<=Wgt_9_489; w_9_490<=Wgt_9_490; w_9_491<=Wgt_9_491; w_9_492<=Wgt_9_492; w_9_493<=Wgt_9_493; w_9_494<=Wgt_9_494; w_9_495<=Wgt_9_495; w_9_496<=Wgt_9_496; w_9_497<=Wgt_9_497; w_9_498<=Wgt_9_498; w_9_499<=Wgt_9_499; w_9_500<=Wgt_9_500; w_9_501<=Wgt_9_501; w_9_502<=Wgt_9_502; w_9_503<=Wgt_9_503; w_9_504<=Wgt_9_504; w_9_505<=Wgt_9_505; w_9_506<=Wgt_9_506; w_9_507<=Wgt_9_507; w_9_508<=Wgt_9_508; w_9_509<=Wgt_9_509; w_9_510<=Wgt_9_510; w_9_511<=Wgt_9_511; w_9_512<=Wgt_9_512; w_9_513<=Wgt_9_513; w_9_514<=Wgt_9_514; w_9_515<=Wgt_9_515; w_9_516<=Wgt_9_516; w_9_517<=Wgt_9_517; w_9_518<=Wgt_9_518; w_9_519<=Wgt_9_519; w_9_520<=Wgt_9_520; w_9_521<=Wgt_9_521; w_9_522<=Wgt_9_522; w_9_523<=Wgt_9_523; w_9_524<=Wgt_9_524; w_9_525<=Wgt_9_525; w_9_526<=Wgt_9_526; w_9_527<=Wgt_9_527; w_9_528<=Wgt_9_528; w_9_529<=Wgt_9_529; w_9_530<=Wgt_9_530; w_9_531<=Wgt_9_531; w_9_532<=Wgt_9_532; w_9_533<=Wgt_9_533; w_9_534<=Wgt_9_534; w_9_535<=Wgt_9_535; w_9_536<=Wgt_9_536; w_9_537<=Wgt_9_537; w_9_538<=Wgt_9_538; w_9_539<=Wgt_9_539; w_9_540<=Wgt_9_540; w_9_541<=Wgt_9_541; w_9_542<=Wgt_9_542; w_9_543<=Wgt_9_543; w_9_544<=Wgt_9_544; w_9_545<=Wgt_9_545; w_9_546<=Wgt_9_546; w_9_547<=Wgt_9_547; w_9_548<=Wgt_9_548; w_9_549<=Wgt_9_549; w_9_550<=Wgt_9_550; w_9_551<=Wgt_9_551; w_9_552<=Wgt_9_552; w_9_553<=Wgt_9_553; w_9_554<=Wgt_9_554; w_9_555<=Wgt_9_555; w_9_556<=Wgt_9_556; w_9_557<=Wgt_9_557; w_9_558<=Wgt_9_558; w_9_559<=Wgt_9_559; w_9_560<=Wgt_9_560; w_9_561<=Wgt_9_561; w_9_562<=Wgt_9_562; w_9_563<=Wgt_9_563; w_9_564<=Wgt_9_564; w_9_565<=Wgt_9_565; w_9_566<=Wgt_9_566; w_9_567<=Wgt_9_567; w_9_568<=Wgt_9_568; w_9_569<=Wgt_9_569; w_9_570<=Wgt_9_570; w_9_571<=Wgt_9_571; w_9_572<=Wgt_9_572; w_9_573<=Wgt_9_573; w_9_574<=Wgt_9_574; w_9_575<=Wgt_9_575; w_9_576<=Wgt_9_576; w_9_577<=Wgt_9_577; w_9_578<=Wgt_9_578; w_9_579<=Wgt_9_579; w_9_580<=Wgt_9_580; w_9_581<=Wgt_9_581; w_9_582<=Wgt_9_582; w_9_583<=Wgt_9_583; w_9_584<=Wgt_9_584; w_9_585<=Wgt_9_585; w_9_586<=Wgt_9_586; w_9_587<=Wgt_9_587; w_9_588<=Wgt_9_588; w_9_589<=Wgt_9_589; w_9_590<=Wgt_9_590; w_9_591<=Wgt_9_591; w_9_592<=Wgt_9_592; w_9_593<=Wgt_9_593; w_9_594<=Wgt_9_594; w_9_595<=Wgt_9_595; w_9_596<=Wgt_9_596; w_9_597<=Wgt_9_597; w_9_598<=Wgt_9_598; w_9_599<=Wgt_9_599; w_9_600<=Wgt_9_600; w_9_601<=Wgt_9_601; w_9_602<=Wgt_9_602; w_9_603<=Wgt_9_603; w_9_604<=Wgt_9_604; w_9_605<=Wgt_9_605; w_9_606<=Wgt_9_606; w_9_607<=Wgt_9_607; w_9_608<=Wgt_9_608; w_9_609<=Wgt_9_609; w_9_610<=Wgt_9_610; w_9_611<=Wgt_9_611; w_9_612<=Wgt_9_612; w_9_613<=Wgt_9_613; w_9_614<=Wgt_9_614; w_9_615<=Wgt_9_615; w_9_616<=Wgt_9_616; w_9_617<=Wgt_9_617; w_9_618<=Wgt_9_618; w_9_619<=Wgt_9_619; w_9_620<=Wgt_9_620; w_9_621<=Wgt_9_621; w_9_622<=Wgt_9_622; w_9_623<=Wgt_9_623; w_9_624<=Wgt_9_624; w_9_625<=Wgt_9_625; w_9_626<=Wgt_9_626; w_9_627<=Wgt_9_627; w_9_628<=Wgt_9_628; w_9_629<=Wgt_9_629; w_9_630<=Wgt_9_630; w_9_631<=Wgt_9_631; w_9_632<=Wgt_9_632; w_9_633<=Wgt_9_633; w_9_634<=Wgt_9_634; w_9_635<=Wgt_9_635; w_9_636<=Wgt_9_636; w_9_637<=Wgt_9_637; w_9_638<=Wgt_9_638; w_9_639<=Wgt_9_639; w_9_640<=Wgt_9_640; w_9_641<=Wgt_9_641; w_9_642<=Wgt_9_642; w_9_643<=Wgt_9_643; w_9_644<=Wgt_9_644; w_9_645<=Wgt_9_645; w_9_646<=Wgt_9_646; w_9_647<=Wgt_9_647; w_9_648<=Wgt_9_648; w_9_649<=Wgt_9_649; w_9_650<=Wgt_9_650; w_9_651<=Wgt_9_651; w_9_652<=Wgt_9_652; w_9_653<=Wgt_9_653; w_9_654<=Wgt_9_654; w_9_655<=Wgt_9_655; w_9_656<=Wgt_9_656; w_9_657<=Wgt_9_657; w_9_658<=Wgt_9_658; w_9_659<=Wgt_9_659; w_9_660<=Wgt_9_660; w_9_661<=Wgt_9_661; w_9_662<=Wgt_9_662; w_9_663<=Wgt_9_663; w_9_664<=Wgt_9_664; w_9_665<=Wgt_9_665; w_9_666<=Wgt_9_666; w_9_667<=Wgt_9_667; w_9_668<=Wgt_9_668; w_9_669<=Wgt_9_669; w_9_670<=Wgt_9_670; w_9_671<=Wgt_9_671; w_9_672<=Wgt_9_672; w_9_673<=Wgt_9_673; w_9_674<=Wgt_9_674; w_9_675<=Wgt_9_675; w_9_676<=Wgt_9_676; w_9_677<=Wgt_9_677; w_9_678<=Wgt_9_678; w_9_679<=Wgt_9_679; w_9_680<=Wgt_9_680; w_9_681<=Wgt_9_681; w_9_682<=Wgt_9_682; w_9_683<=Wgt_9_683; w_9_684<=Wgt_9_684; w_9_685<=Wgt_9_685; w_9_686<=Wgt_9_686; w_9_687<=Wgt_9_687; w_9_688<=Wgt_9_688; w_9_689<=Wgt_9_689; w_9_690<=Wgt_9_690; w_9_691<=Wgt_9_691; w_9_692<=Wgt_9_692; w_9_693<=Wgt_9_693; w_9_694<=Wgt_9_694; w_9_695<=Wgt_9_695; w_9_696<=Wgt_9_696; w_9_697<=Wgt_9_697; w_9_698<=Wgt_9_698; w_9_699<=Wgt_9_699; w_9_700<=Wgt_9_700; w_9_701<=Wgt_9_701; w_9_702<=Wgt_9_702; w_9_703<=Wgt_9_703; w_9_704<=Wgt_9_704; w_9_705<=Wgt_9_705; w_9_706<=Wgt_9_706; w_9_707<=Wgt_9_707; w_9_708<=Wgt_9_708; w_9_709<=Wgt_9_709; w_9_710<=Wgt_9_710; w_9_711<=Wgt_9_711; w_9_712<=Wgt_9_712; w_9_713<=Wgt_9_713; w_9_714<=Wgt_9_714; w_9_715<=Wgt_9_715; w_9_716<=Wgt_9_716; w_9_717<=Wgt_9_717; w_9_718<=Wgt_9_718; w_9_719<=Wgt_9_719; w_9_720<=Wgt_9_720; w_9_721<=Wgt_9_721; w_9_722<=Wgt_9_722; w_9_723<=Wgt_9_723; w_9_724<=Wgt_9_724; w_9_725<=Wgt_9_725; w_9_726<=Wgt_9_726; w_9_727<=Wgt_9_727; w_9_728<=Wgt_9_728; w_9_729<=Wgt_9_729; w_9_730<=Wgt_9_730; w_9_731<=Wgt_9_731; w_9_732<=Wgt_9_732; w_9_733<=Wgt_9_733; w_9_734<=Wgt_9_734; w_9_735<=Wgt_9_735; w_9_736<=Wgt_9_736; w_9_737<=Wgt_9_737; w_9_738<=Wgt_9_738; w_9_739<=Wgt_9_739; w_9_740<=Wgt_9_740; w_9_741<=Wgt_9_741; w_9_742<=Wgt_9_742; w_9_743<=Wgt_9_743; w_9_744<=Wgt_9_744; w_9_745<=Wgt_9_745; w_9_746<=Wgt_9_746; w_9_747<=Wgt_9_747; w_9_748<=Wgt_9_748; w_9_749<=Wgt_9_749; w_9_750<=Wgt_9_750; w_9_751<=Wgt_9_751; w_9_752<=Wgt_9_752; w_9_753<=Wgt_9_753; w_9_754<=Wgt_9_754; w_9_755<=Wgt_9_755; w_9_756<=Wgt_9_756; w_9_757<=Wgt_9_757; w_9_758<=Wgt_9_758; w_9_759<=Wgt_9_759; w_9_760<=Wgt_9_760; w_9_761<=Wgt_9_761; w_9_762<=Wgt_9_762; w_9_763<=Wgt_9_763; w_9_764<=Wgt_9_764; w_9_765<=Wgt_9_765; w_9_766<=Wgt_9_766; w_9_767<=Wgt_9_767; w_9_768<=Wgt_9_768; w_9_769<=Wgt_9_769; w_9_770<=Wgt_9_770; w_9_771<=Wgt_9_771; w_9_772<=Wgt_9_772; w_9_773<=Wgt_9_773; w_9_774<=Wgt_9_774; w_9_775<=Wgt_9_775; w_9_776<=Wgt_9_776; w_9_777<=Wgt_9_777; w_9_778<=Wgt_9_778; w_9_779<=Wgt_9_779; w_9_780<=Wgt_9_780; w_9_781<=Wgt_9_781; w_9_782<=Wgt_9_782; w_9_783<=Wgt_9_783; w_9_784<=Wgt_9_784; 
					//select<=select+1; 
				end
			else
			begin
			end
		end
end		
//input to register
always @(posedge clk or negedge GlobalReset) begin
	if (GlobalReset == 1'b0)
		begin
			select <= 0;
		end
	else

		begin
		
			case(select)
			//input everything to regist during 1st clk
				8'd0: 	if(Input_Valid)
						begin
						//input all pixel value
						select<=select+1; 
						end
						else
						begin
						select<=8'd0;
						end
				8'd1:
					begin
						wr0<=w_0_0; wr1<=w_0_1; wr2<=w_0_2; wr3<=w_0_3; wr4<=w_0_4; wr5<=w_0_5; wr6<=w_0_6; wr7<=w_0_7; wr8<=w_0_8; wr9<=w_0_9; wr10<=w_0_10; wr11<=w_0_11; wr12<=w_0_12; wr13<=w_0_13; wr14<=w_0_14; wr15<=w_0_15; wr16<=w_0_16; wr17<=w_0_17; wr18<=w_0_18; wr19<=w_0_19; wr20<=w_0_20; wr21<=w_0_21; wr22<=w_0_22; wr23<=w_0_23; wr24<=w_0_24; wr25<=w_0_25; wr26<=w_0_26; wr27<=w_0_27; wr28<=w_0_28; wr29<=w_0_29; wr30<=w_0_30; wr31<=w_0_31; wr32<=w_0_32; wr33<=w_0_33; wr34<=w_0_34; wr35<=w_0_35; wr36<=w_0_36; wr37<=w_0_37; wr38<=w_0_38; wr39<=w_0_39; wr40<=w_0_40; wr41<=w_0_41; wr42<=w_0_42; wr43<=w_0_43; wr44<=w_0_44; wr45<=w_0_45; wr46<=w_0_46; wr47<=w_0_47; wr48<=w_0_48; wr49<=w_0_49; wr50<=w_0_50; wr51<=w_0_51; wr52<=w_0_52; wr53<=w_0_53; wr54<=w_0_54; wr55<=w_0_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd2:
					begin
						wr0<=w_0_56; wr1<=w_0_57; wr2<=w_0_58; wr3<=w_0_59; wr4<=w_0_60; wr5<=w_0_61; wr6<=w_0_62; wr7<=w_0_63; wr8<=w_0_64; wr9<=w_0_65; wr10<=w_0_66; wr11<=w_0_67; wr12<=w_0_68; wr13<=w_0_69; wr14<=w_0_70; wr15<=w_0_71; wr16<=w_0_72; wr17<=w_0_73; wr18<=w_0_74; wr19<=w_0_75; wr20<=w_0_76; wr21<=w_0_77; wr22<=w_0_78; wr23<=w_0_79; wr24<=w_0_80; wr25<=w_0_81; wr26<=w_0_82; wr27<=w_0_83; wr28<=w_0_84; wr29<=w_0_85; wr30<=w_0_86; wr31<=w_0_87; wr32<=w_0_88; wr33<=w_0_89; wr34<=w_0_90; wr35<=w_0_91; wr36<=w_0_92; wr37<=w_0_93; wr38<=w_0_94; wr39<=w_0_95; wr40<=w_0_96; wr41<=w_0_97; wr42<=w_0_98; wr43<=w_0_99; wr44<=w_0_100; wr45<=w_0_101; wr46<=w_0_102; wr47<=w_0_103; wr48<=w_0_104; wr49<=w_0_105; wr50<=w_0_106; wr51<=w_0_107; wr52<=w_0_108; wr53<=w_0_109; wr54<=w_0_110; wr55<=w_0_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd3:
					begin
						wr0<=w_0_112; wr1<=w_0_113; wr2<=w_0_114; wr3<=w_0_115; wr4<=w_0_116; wr5<=w_0_117; wr6<=w_0_118; wr7<=w_0_119; wr8<=w_0_120; wr9<=w_0_121; wr10<=w_0_122; wr11<=w_0_123; wr12<=w_0_124; wr13<=w_0_125; wr14<=w_0_126; wr15<=w_0_127; wr16<=w_0_128; wr17<=w_0_129; wr18<=w_0_130; wr19<=w_0_131; wr20<=w_0_132; wr21<=w_0_133; wr22<=w_0_134; wr23<=w_0_135; wr24<=w_0_136; wr25<=w_0_137; wr26<=w_0_138; wr27<=w_0_139; wr28<=w_0_140; wr29<=w_0_141; wr30<=w_0_142; wr31<=w_0_143; wr32<=w_0_144; wr33<=w_0_145; wr34<=w_0_146; wr35<=w_0_147; wr36<=w_0_148; wr37<=w_0_149; wr38<=w_0_150; wr39<=w_0_151; wr40<=w_0_152; wr41<=w_0_153; wr42<=w_0_154; wr43<=w_0_155; wr44<=w_0_156; wr45<=w_0_157; wr46<=w_0_158; wr47<=w_0_159; wr48<=w_0_160; wr49<=w_0_161; wr50<=w_0_162; wr51<=w_0_163; wr52<=w_0_164; wr53<=w_0_165; wr54<=w_0_166; wr55<=w_0_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd4:
					begin
						wr0<=w_0_168; wr1<=w_0_169; wr2<=w_0_170; wr3<=w_0_171; wr4<=w_0_172; wr5<=w_0_173; wr6<=w_0_174; wr7<=w_0_175; wr8<=w_0_176; wr9<=w_0_177; wr10<=w_0_178; wr11<=w_0_179; wr12<=w_0_180; wr13<=w_0_181; wr14<=w_0_182; wr15<=w_0_183; wr16<=w_0_184; wr17<=w_0_185; wr18<=w_0_186; wr19<=w_0_187; wr20<=w_0_188; wr21<=w_0_189; wr22<=w_0_190; wr23<=w_0_191; wr24<=w_0_192; wr25<=w_0_193; wr26<=w_0_194; wr27<=w_0_195; wr28<=w_0_196; wr29<=w_0_197; wr30<=w_0_198; wr31<=w_0_199; wr32<=w_0_200; wr33<=w_0_201; wr34<=w_0_202; wr35<=w_0_203; wr36<=w_0_204; wr37<=w_0_205; wr38<=w_0_206; wr39<=w_0_207; wr40<=w_0_208; wr41<=w_0_209; wr42<=w_0_210; wr43<=w_0_211; wr44<=w_0_212; wr45<=w_0_213; wr46<=w_0_214; wr47<=w_0_215; wr48<=w_0_216; wr49<=w_0_217; wr50<=w_0_218; wr51<=w_0_219; wr52<=w_0_220; wr53<=w_0_221; wr54<=w_0_222; wr55<=w_0_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd5:
					begin
						wr0<=w_0_224; wr1<=w_0_225; wr2<=w_0_226; wr3<=w_0_227; wr4<=w_0_228; wr5<=w_0_229; wr6<=w_0_230; wr7<=w_0_231; wr8<=w_0_232; wr9<=w_0_233; wr10<=w_0_234; wr11<=w_0_235; wr12<=w_0_236; wr13<=w_0_237; wr14<=w_0_238; wr15<=w_0_239; wr16<=w_0_240; wr17<=w_0_241; wr18<=w_0_242; wr19<=w_0_243; wr20<=w_0_244; wr21<=w_0_245; wr22<=w_0_246; wr23<=w_0_247; wr24<=w_0_248; wr25<=w_0_249; wr26<=w_0_250; wr27<=w_0_251; wr28<=w_0_252; wr29<=w_0_253; wr30<=w_0_254; wr31<=w_0_255; wr32<=w_0_256; wr33<=w_0_257; wr34<=w_0_258; wr35<=w_0_259; wr36<=w_0_260; wr37<=w_0_261; wr38<=w_0_262; wr39<=w_0_263; wr40<=w_0_264; wr41<=w_0_265; wr42<=w_0_266; wr43<=w_0_267; wr44<=w_0_268; wr45<=w_0_269; wr46<=w_0_270; wr47<=w_0_271; wr48<=w_0_272; wr49<=w_0_273; wr50<=w_0_274; wr51<=w_0_275; wr52<=w_0_276; wr53<=w_0_277; wr54<=w_0_278; wr55<=w_0_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd6:
					begin
						wr0<=w_0_280; wr1<=w_0_281; wr2<=w_0_282; wr3<=w_0_283; wr4<=w_0_284; wr5<=w_0_285; wr6<=w_0_286; wr7<=w_0_287; wr8<=w_0_288; wr9<=w_0_289; wr10<=w_0_290; wr11<=w_0_291; wr12<=w_0_292; wr13<=w_0_293; wr14<=w_0_294; wr15<=w_0_295; wr16<=w_0_296; wr17<=w_0_297; wr18<=w_0_298; wr19<=w_0_299; wr20<=w_0_300; wr21<=w_0_301; wr22<=w_0_302; wr23<=w_0_303; wr24<=w_0_304; wr25<=w_0_305; wr26<=w_0_306; wr27<=w_0_307; wr28<=w_0_308; wr29<=w_0_309; wr30<=w_0_310; wr31<=w_0_311; wr32<=w_0_312; wr33<=w_0_313; wr34<=w_0_314; wr35<=w_0_315; wr36<=w_0_316; wr37<=w_0_317; wr38<=w_0_318; wr39<=w_0_319; wr40<=w_0_320; wr41<=w_0_321; wr42<=w_0_322; wr43<=w_0_323; wr44<=w_0_324; wr45<=w_0_325; wr46<=w_0_326; wr47<=w_0_327; wr48<=w_0_328; wr49<=w_0_329; wr50<=w_0_330; wr51<=w_0_331; wr52<=w_0_332; wr53<=w_0_333; wr54<=w_0_334; wr55<=w_0_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd7:
					begin
						wr0<=w_0_336; wr1<=w_0_337; wr2<=w_0_338; wr3<=w_0_339; wr4<=w_0_340; wr5<=w_0_341; wr6<=w_0_342; wr7<=w_0_343; wr8<=w_0_344; wr9<=w_0_345; wr10<=w_0_346; wr11<=w_0_347; wr12<=w_0_348; wr13<=w_0_349; wr14<=w_0_350; wr15<=w_0_351; wr16<=w_0_352; wr17<=w_0_353; wr18<=w_0_354; wr19<=w_0_355; wr20<=w_0_356; wr21<=w_0_357; wr22<=w_0_358; wr23<=w_0_359; wr24<=w_0_360; wr25<=w_0_361; wr26<=w_0_362; wr27<=w_0_363; wr28<=w_0_364; wr29<=w_0_365; wr30<=w_0_366; wr31<=w_0_367; wr32<=w_0_368; wr33<=w_0_369; wr34<=w_0_370; wr35<=w_0_371; wr36<=w_0_372; wr37<=w_0_373; wr38<=w_0_374; wr39<=w_0_375; wr40<=w_0_376; wr41<=w_0_377; wr42<=w_0_378; wr43<=w_0_379; wr44<=w_0_380; wr45<=w_0_381; wr46<=w_0_382; wr47<=w_0_383; wr48<=w_0_384; wr49<=w_0_385; wr50<=w_0_386; wr51<=w_0_387; wr52<=w_0_388; wr53<=w_0_389; wr54<=w_0_390; wr55<=w_0_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd8:
					begin
						wr0<=w_0_392; wr1<=w_0_393; wr2<=w_0_394; wr3<=w_0_395; wr4<=w_0_396; wr5<=w_0_397; wr6<=w_0_398; wr7<=w_0_399; wr8<=w_0_400; wr9<=w_0_401; wr10<=w_0_402; wr11<=w_0_403; wr12<=w_0_404; wr13<=w_0_405; wr14<=w_0_406; wr15<=w_0_407; wr16<=w_0_408; wr17<=w_0_409; wr18<=w_0_410; wr19<=w_0_411; wr20<=w_0_412; wr21<=w_0_413; wr22<=w_0_414; wr23<=w_0_415; wr24<=w_0_416; wr25<=w_0_417; wr26<=w_0_418; wr27<=w_0_419; wr28<=w_0_420; wr29<=w_0_421; wr30<=w_0_422; wr31<=w_0_423; wr32<=w_0_424; wr33<=w_0_425; wr34<=w_0_426; wr35<=w_0_427; wr36<=w_0_428; wr37<=w_0_429; wr38<=w_0_430; wr39<=w_0_431; wr40<=w_0_432; wr41<=w_0_433; wr42<=w_0_434; wr43<=w_0_435; wr44<=w_0_436; wr45<=w_0_437; wr46<=w_0_438; wr47<=w_0_439; wr48<=w_0_440; wr49<=w_0_441; wr50<=w_0_442; wr51<=w_0_443; wr52<=w_0_444; wr53<=w_0_445; wr54<=w_0_446; wr55<=w_0_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd9:
					begin
						wr0<=w_0_448; wr1<=w_0_449; wr2<=w_0_450; wr3<=w_0_451; wr4<=w_0_452; wr5<=w_0_453; wr6<=w_0_454; wr7<=w_0_455; wr8<=w_0_456; wr9<=w_0_457; wr10<=w_0_458; wr11<=w_0_459; wr12<=w_0_460; wr13<=w_0_461; wr14<=w_0_462; wr15<=w_0_463; wr16<=w_0_464; wr17<=w_0_465; wr18<=w_0_466; wr19<=w_0_467; wr20<=w_0_468; wr21<=w_0_469; wr22<=w_0_470; wr23<=w_0_471; wr24<=w_0_472; wr25<=w_0_473; wr26<=w_0_474; wr27<=w_0_475; wr28<=w_0_476; wr29<=w_0_477; wr30<=w_0_478; wr31<=w_0_479; wr32<=w_0_480; wr33<=w_0_481; wr34<=w_0_482; wr35<=w_0_483; wr36<=w_0_484; wr37<=w_0_485; wr38<=w_0_486; wr39<=w_0_487; wr40<=w_0_488; wr41<=w_0_489; wr42<=w_0_490; wr43<=w_0_491; wr44<=w_0_492; wr45<=w_0_493; wr46<=w_0_494; wr47<=w_0_495; wr48<=w_0_496; wr49<=w_0_497; wr50<=w_0_498; wr51<=w_0_499; wr52<=w_0_500; wr53<=w_0_501; wr54<=w_0_502; wr55<=w_0_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd10:
					begin
						wr0<=w_0_504; wr1<=w_0_505; wr2<=w_0_506; wr3<=w_0_507; wr4<=w_0_508; wr5<=w_0_509; wr6<=w_0_510; wr7<=w_0_511; wr8<=w_0_512; wr9<=w_0_513; wr10<=w_0_514; wr11<=w_0_515; wr12<=w_0_516; wr13<=w_0_517; wr14<=w_0_518; wr15<=w_0_519; wr16<=w_0_520; wr17<=w_0_521; wr18<=w_0_522; wr19<=w_0_523; wr20<=w_0_524; wr21<=w_0_525; wr22<=w_0_526; wr23<=w_0_527; wr24<=w_0_528; wr25<=w_0_529; wr26<=w_0_530; wr27<=w_0_531; wr28<=w_0_532; wr29<=w_0_533; wr30<=w_0_534; wr31<=w_0_535; wr32<=w_0_536; wr33<=w_0_537; wr34<=w_0_538; wr35<=w_0_539; wr36<=w_0_540; wr37<=w_0_541; wr38<=w_0_542; wr39<=w_0_543; wr40<=w_0_544; wr41<=w_0_545; wr42<=w_0_546; wr43<=w_0_547; wr44<=w_0_548; wr45<=w_0_549; wr46<=w_0_550; wr47<=w_0_551; wr48<=w_0_552; wr49<=w_0_553; wr50<=w_0_554; wr51<=w_0_555; wr52<=w_0_556; wr53<=w_0_557; wr54<=w_0_558; wr55<=w_0_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd11:
					begin
						wr0<=w_0_560; wr1<=w_0_561; wr2<=w_0_562; wr3<=w_0_563; wr4<=w_0_564; wr5<=w_0_565; wr6<=w_0_566; wr7<=w_0_567; wr8<=w_0_568; wr9<=w_0_569; wr10<=w_0_570; wr11<=w_0_571; wr12<=w_0_572; wr13<=w_0_573; wr14<=w_0_574; wr15<=w_0_575; wr16<=w_0_576; wr17<=w_0_577; wr18<=w_0_578; wr19<=w_0_579; wr20<=w_0_580; wr21<=w_0_581; wr22<=w_0_582; wr23<=w_0_583; wr24<=w_0_584; wr25<=w_0_585; wr26<=w_0_586; wr27<=w_0_587; wr28<=w_0_588; wr29<=w_0_589; wr30<=w_0_590; wr31<=w_0_591; wr32<=w_0_592; wr33<=w_0_593; wr34<=w_0_594; wr35<=w_0_595; wr36<=w_0_596; wr37<=w_0_597; wr38<=w_0_598; wr39<=w_0_599; wr40<=w_0_600; wr41<=w_0_601; wr42<=w_0_602; wr43<=w_0_603; wr44<=w_0_604; wr45<=w_0_605; wr46<=w_0_606; wr47<=w_0_607; wr48<=w_0_608; wr49<=w_0_609; wr50<=w_0_610; wr51<=w_0_611; wr52<=w_0_612; wr53<=w_0_613; wr54<=w_0_614; wr55<=w_0_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd12:
					begin
						wr0<=w_0_616; wr1<=w_0_617; wr2<=w_0_618; wr3<=w_0_619; wr4<=w_0_620; wr5<=w_0_621; wr6<=w_0_622; wr7<=w_0_623; wr8<=w_0_624; wr9<=w_0_625; wr10<=w_0_626; wr11<=w_0_627; wr12<=w_0_628; wr13<=w_0_629; wr14<=w_0_630; wr15<=w_0_631; wr16<=w_0_632; wr17<=w_0_633; wr18<=w_0_634; wr19<=w_0_635; wr20<=w_0_636; wr21<=w_0_637; wr22<=w_0_638; wr23<=w_0_639; wr24<=w_0_640; wr25<=w_0_641; wr26<=w_0_642; wr27<=w_0_643; wr28<=w_0_644; wr29<=w_0_645; wr30<=w_0_646; wr31<=w_0_647; wr32<=w_0_648; wr33<=w_0_649; wr34<=w_0_650; wr35<=w_0_651; wr36<=w_0_652; wr37<=w_0_653; wr38<=w_0_654; wr39<=w_0_655; wr40<=w_0_656; wr41<=w_0_657; wr42<=w_0_658; wr43<=w_0_659; wr44<=w_0_660; wr45<=w_0_661; wr46<=w_0_662; wr47<=w_0_663; wr48<=w_0_664; wr49<=w_0_665; wr50<=w_0_666; wr51<=w_0_667; wr52<=w_0_668; wr53<=w_0_669; wr54<=w_0_670; wr55<=w_0_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd13:
					begin
						wr0<=w_0_672; wr1<=w_0_673; wr2<=w_0_674; wr3<=w_0_675; wr4<=w_0_676; wr5<=w_0_677; wr6<=w_0_678; wr7<=w_0_679; wr8<=w_0_680; wr9<=w_0_681; wr10<=w_0_682; wr11<=w_0_683; wr12<=w_0_684; wr13<=w_0_685; wr14<=w_0_686; wr15<=w_0_687; wr16<=w_0_688; wr17<=w_0_689; wr18<=w_0_690; wr19<=w_0_691; wr20<=w_0_692; wr21<=w_0_693; wr22<=w_0_694; wr23<=w_0_695; wr24<=w_0_696; wr25<=w_0_697; wr26<=w_0_698; wr27<=w_0_699; wr28<=w_0_700; wr29<=w_0_701; wr30<=w_0_702; wr31<=w_0_703; wr32<=w_0_704; wr33<=w_0_705; wr34<=w_0_706; wr35<=w_0_707; wr36<=w_0_708; wr37<=w_0_709; wr38<=w_0_710; wr39<=w_0_711; wr40<=w_0_712; wr41<=w_0_713; wr42<=w_0_714; wr43<=w_0_715; wr44<=w_0_716; wr45<=w_0_717; wr46<=w_0_718; wr47<=w_0_719; wr48<=w_0_720; wr49<=w_0_721; wr50<=w_0_722; wr51<=w_0_723; wr52<=w_0_724; wr53<=w_0_725; wr54<=w_0_726; wr55<=w_0_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd14:
					begin
						wr0<=w_0_728; wr1<=w_0_729; wr2<=w_0_730; wr3<=w_0_731; wr4<=w_0_732; wr5<=w_0_733; wr6<=w_0_734; wr7<=w_0_735; wr8<=w_0_736; wr9<=w_0_737; wr10<=w_0_738; wr11<=w_0_739; wr12<=w_0_740; wr13<=w_0_741; wr14<=w_0_742; wr15<=w_0_743; wr16<=w_0_744; wr17<=w_0_745; wr18<=w_0_746; wr19<=w_0_747; wr20<=w_0_748; wr21<=w_0_749; wr22<=w_0_750; wr23<=w_0_751; wr24<=w_0_752; wr25<=w_0_753; wr26<=w_0_754; wr27<=w_0_755; wr28<=w_0_756; wr29<=w_0_757; wr30<=w_0_758; wr31<=w_0_759; wr32<=w_0_760; wr33<=w_0_761; wr34<=w_0_762; wr35<=w_0_763; wr36<=w_0_764; wr37<=w_0_765; wr38<=w_0_766; wr39<=w_0_767; wr40<=w_0_768; wr41<=w_0_769; wr42<=w_0_770; wr43<=w_0_771; wr44<=w_0_772; wr45<=w_0_773; wr46<=w_0_774; wr47<=w_0_775; wr48<=w_0_776; wr49<=w_0_777; wr50<=w_0_778; wr51<=w_0_779; wr52<=w_0_780; wr53<=w_0_781; wr54<=w_0_782; wr55<=w_0_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd15:
					begin
						bias_p<=px_784;
						bias_w<=w_0_784;
						select<=select+1;
					end
				8'd16:
					begin
						wr0<=w_1_0; wr1<=w_1_1; wr2<=w_1_2; wr3<=w_1_3; wr4<=w_1_4; wr5<=w_1_5; wr6<=w_1_6; wr7<=w_1_7; wr8<=w_1_8; wr9<=w_1_9; wr10<=w_1_10; wr11<=w_1_11; wr12<=w_1_12; wr13<=w_1_13; wr14<=w_1_14; wr15<=w_1_15; wr16<=w_1_16; wr17<=w_1_17; wr18<=w_1_18; wr19<=w_1_19; wr20<=w_1_20; wr21<=w_1_21; wr22<=w_1_22; wr23<=w_1_23; wr24<=w_1_24; wr25<=w_1_25; wr26<=w_1_26; wr27<=w_1_27; wr28<=w_1_28; wr29<=w_1_29; wr30<=w_1_30; wr31<=w_1_31; wr32<=w_1_32; wr33<=w_1_33; wr34<=w_1_34; wr35<=w_1_35; wr36<=w_1_36; wr37<=w_1_37; wr38<=w_1_38; wr39<=w_1_39; wr40<=w_1_40; wr41<=w_1_41; wr42<=w_1_42; wr43<=w_1_43; wr44<=w_1_44; wr45<=w_1_45; wr46<=w_1_46; wr47<=w_1_47; wr48<=w_1_48; wr49<=w_1_49; wr50<=w_1_50; wr51<=w_1_51; wr52<=w_1_52; wr53<=w_1_53; wr54<=w_1_54; wr55<=w_1_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd17:
					begin
						wr0<=w_1_56; wr1<=w_1_57; wr2<=w_1_58; wr3<=w_1_59; wr4<=w_1_60; wr5<=w_1_61; wr6<=w_1_62; wr7<=w_1_63; wr8<=w_1_64; wr9<=w_1_65; wr10<=w_1_66; wr11<=w_1_67; wr12<=w_1_68; wr13<=w_1_69; wr14<=w_1_70; wr15<=w_1_71; wr16<=w_1_72; wr17<=w_1_73; wr18<=w_1_74; wr19<=w_1_75; wr20<=w_1_76; wr21<=w_1_77; wr22<=w_1_78; wr23<=w_1_79; wr24<=w_1_80; wr25<=w_1_81; wr26<=w_1_82; wr27<=w_1_83; wr28<=w_1_84; wr29<=w_1_85; wr30<=w_1_86; wr31<=w_1_87; wr32<=w_1_88; wr33<=w_1_89; wr34<=w_1_90; wr35<=w_1_91; wr36<=w_1_92; wr37<=w_1_93; wr38<=w_1_94; wr39<=w_1_95; wr40<=w_1_96; wr41<=w_1_97; wr42<=w_1_98; wr43<=w_1_99; wr44<=w_1_100; wr45<=w_1_101; wr46<=w_1_102; wr47<=w_1_103; wr48<=w_1_104; wr49<=w_1_105; wr50<=w_1_106; wr51<=w_1_107; wr52<=w_1_108; wr53<=w_1_109; wr54<=w_1_110; wr55<=w_1_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd18:
					begin
						wr0<=w_1_112; wr1<=w_1_113; wr2<=w_1_114; wr3<=w_1_115; wr4<=w_1_116; wr5<=w_1_117; wr6<=w_1_118; wr7<=w_1_119; wr8<=w_1_120; wr9<=w_1_121; wr10<=w_1_122; wr11<=w_1_123; wr12<=w_1_124; wr13<=w_1_125; wr14<=w_1_126; wr15<=w_1_127; wr16<=w_1_128; wr17<=w_1_129; wr18<=w_1_130; wr19<=w_1_131; wr20<=w_1_132; wr21<=w_1_133; wr22<=w_1_134; wr23<=w_1_135; wr24<=w_1_136; wr25<=w_1_137; wr26<=w_1_138; wr27<=w_1_139; wr28<=w_1_140; wr29<=w_1_141; wr30<=w_1_142; wr31<=w_1_143; wr32<=w_1_144; wr33<=w_1_145; wr34<=w_1_146; wr35<=w_1_147; wr36<=w_1_148; wr37<=w_1_149; wr38<=w_1_150; wr39<=w_1_151; wr40<=w_1_152; wr41<=w_1_153; wr42<=w_1_154; wr43<=w_1_155; wr44<=w_1_156; wr45<=w_1_157; wr46<=w_1_158; wr47<=w_1_159; wr48<=w_1_160; wr49<=w_1_161; wr50<=w_1_162; wr51<=w_1_163; wr52<=w_1_164; wr53<=w_1_165; wr54<=w_1_166; wr55<=w_1_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd19:
					begin
						wr0<=w_1_168; wr1<=w_1_169; wr2<=w_1_170; wr3<=w_1_171; wr4<=w_1_172; wr5<=w_1_173; wr6<=w_1_174; wr7<=w_1_175; wr8<=w_1_176; wr9<=w_1_177; wr10<=w_1_178; wr11<=w_1_179; wr12<=w_1_180; wr13<=w_1_181; wr14<=w_1_182; wr15<=w_1_183; wr16<=w_1_184; wr17<=w_1_185; wr18<=w_1_186; wr19<=w_1_187; wr20<=w_1_188; wr21<=w_1_189; wr22<=w_1_190; wr23<=w_1_191; wr24<=w_1_192; wr25<=w_1_193; wr26<=w_1_194; wr27<=w_1_195; wr28<=w_1_196; wr29<=w_1_197; wr30<=w_1_198; wr31<=w_1_199; wr32<=w_1_200; wr33<=w_1_201; wr34<=w_1_202; wr35<=w_1_203; wr36<=w_1_204; wr37<=w_1_205; wr38<=w_1_206; wr39<=w_1_207; wr40<=w_1_208; wr41<=w_1_209; wr42<=w_1_210; wr43<=w_1_211; wr44<=w_1_212; wr45<=w_1_213; wr46<=w_1_214; wr47<=w_1_215; wr48<=w_1_216; wr49<=w_1_217; wr50<=w_1_218; wr51<=w_1_219; wr52<=w_1_220; wr53<=w_1_221; wr54<=w_1_222; wr55<=w_1_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd20:
					begin
						wr0<=w_1_224; wr1<=w_1_225; wr2<=w_1_226; wr3<=w_1_227; wr4<=w_1_228; wr5<=w_1_229; wr6<=w_1_230; wr7<=w_1_231; wr8<=w_1_232; wr9<=w_1_233; wr10<=w_1_234; wr11<=w_1_235; wr12<=w_1_236; wr13<=w_1_237; wr14<=w_1_238; wr15<=w_1_239; wr16<=w_1_240; wr17<=w_1_241; wr18<=w_1_242; wr19<=w_1_243; wr20<=w_1_244; wr21<=w_1_245; wr22<=w_1_246; wr23<=w_1_247; wr24<=w_1_248; wr25<=w_1_249; wr26<=w_1_250; wr27<=w_1_251; wr28<=w_1_252; wr29<=w_1_253; wr30<=w_1_254; wr31<=w_1_255; wr32<=w_1_256; wr33<=w_1_257; wr34<=w_1_258; wr35<=w_1_259; wr36<=w_1_260; wr37<=w_1_261; wr38<=w_1_262; wr39<=w_1_263; wr40<=w_1_264; wr41<=w_1_265; wr42<=w_1_266; wr43<=w_1_267; wr44<=w_1_268; wr45<=w_1_269; wr46<=w_1_270; wr47<=w_1_271; wr48<=w_1_272; wr49<=w_1_273; wr50<=w_1_274; wr51<=w_1_275; wr52<=w_1_276; wr53<=w_1_277; wr54<=w_1_278; wr55<=w_1_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd21:
					begin
						wr0<=w_1_280; wr1<=w_1_281; wr2<=w_1_282; wr3<=w_1_283; wr4<=w_1_284; wr5<=w_1_285; wr6<=w_1_286; wr7<=w_1_287; wr8<=w_1_288; wr9<=w_1_289; wr10<=w_1_290; wr11<=w_1_291; wr12<=w_1_292; wr13<=w_1_293; wr14<=w_1_294; wr15<=w_1_295; wr16<=w_1_296; wr17<=w_1_297; wr18<=w_1_298; wr19<=w_1_299; wr20<=w_1_300; wr21<=w_1_301; wr22<=w_1_302; wr23<=w_1_303; wr24<=w_1_304; wr25<=w_1_305; wr26<=w_1_306; wr27<=w_1_307; wr28<=w_1_308; wr29<=w_1_309; wr30<=w_1_310; wr31<=w_1_311; wr32<=w_1_312; wr33<=w_1_313; wr34<=w_1_314; wr35<=w_1_315; wr36<=w_1_316; wr37<=w_1_317; wr38<=w_1_318; wr39<=w_1_319; wr40<=w_1_320; wr41<=w_1_321; wr42<=w_1_322; wr43<=w_1_323; wr44<=w_1_324; wr45<=w_1_325; wr46<=w_1_326; wr47<=w_1_327; wr48<=w_1_328; wr49<=w_1_329; wr50<=w_1_330; wr51<=w_1_331; wr52<=w_1_332; wr53<=w_1_333; wr54<=w_1_334; wr55<=w_1_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd22:
					begin
						wr0<=w_1_336; wr1<=w_1_337; wr2<=w_1_338; wr3<=w_1_339; wr4<=w_1_340; wr5<=w_1_341; wr6<=w_1_342; wr7<=w_1_343; wr8<=w_1_344; wr9<=w_1_345; wr10<=w_1_346; wr11<=w_1_347; wr12<=w_1_348; wr13<=w_1_349; wr14<=w_1_350; wr15<=w_1_351; wr16<=w_1_352; wr17<=w_1_353; wr18<=w_1_354; wr19<=w_1_355; wr20<=w_1_356; wr21<=w_1_357; wr22<=w_1_358; wr23<=w_1_359; wr24<=w_1_360; wr25<=w_1_361; wr26<=w_1_362; wr27<=w_1_363; wr28<=w_1_364; wr29<=w_1_365; wr30<=w_1_366; wr31<=w_1_367; wr32<=w_1_368; wr33<=w_1_369; wr34<=w_1_370; wr35<=w_1_371; wr36<=w_1_372; wr37<=w_1_373; wr38<=w_1_374; wr39<=w_1_375; wr40<=w_1_376; wr41<=w_1_377; wr42<=w_1_378; wr43<=w_1_379; wr44<=w_1_380; wr45<=w_1_381; wr46<=w_1_382; wr47<=w_1_383; wr48<=w_1_384; wr49<=w_1_385; wr50<=w_1_386; wr51<=w_1_387; wr52<=w_1_388; wr53<=w_1_389; wr54<=w_1_390; wr55<=w_1_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd23:
					begin
						wr0<=w_1_392; wr1<=w_1_393; wr2<=w_1_394; wr3<=w_1_395; wr4<=w_1_396; wr5<=w_1_397; wr6<=w_1_398; wr7<=w_1_399; wr8<=w_1_400; wr9<=w_1_401; wr10<=w_1_402; wr11<=w_1_403; wr12<=w_1_404; wr13<=w_1_405; wr14<=w_1_406; wr15<=w_1_407; wr16<=w_1_408; wr17<=w_1_409; wr18<=w_1_410; wr19<=w_1_411; wr20<=w_1_412; wr21<=w_1_413; wr22<=w_1_414; wr23<=w_1_415; wr24<=w_1_416; wr25<=w_1_417; wr26<=w_1_418; wr27<=w_1_419; wr28<=w_1_420; wr29<=w_1_421; wr30<=w_1_422; wr31<=w_1_423; wr32<=w_1_424; wr33<=w_1_425; wr34<=w_1_426; wr35<=w_1_427; wr36<=w_1_428; wr37<=w_1_429; wr38<=w_1_430; wr39<=w_1_431; wr40<=w_1_432; wr41<=w_1_433; wr42<=w_1_434; wr43<=w_1_435; wr44<=w_1_436; wr45<=w_1_437; wr46<=w_1_438; wr47<=w_1_439; wr48<=w_1_440; wr49<=w_1_441; wr50<=w_1_442; wr51<=w_1_443; wr52<=w_1_444; wr53<=w_1_445; wr54<=w_1_446; wr55<=w_1_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd24:
					begin
						wr0<=w_1_448; wr1<=w_1_449; wr2<=w_1_450; wr3<=w_1_451; wr4<=w_1_452; wr5<=w_1_453; wr6<=w_1_454; wr7<=w_1_455; wr8<=w_1_456; wr9<=w_1_457; wr10<=w_1_458; wr11<=w_1_459; wr12<=w_1_460; wr13<=w_1_461; wr14<=w_1_462; wr15<=w_1_463; wr16<=w_1_464; wr17<=w_1_465; wr18<=w_1_466; wr19<=w_1_467; wr20<=w_1_468; wr21<=w_1_469; wr22<=w_1_470; wr23<=w_1_471; wr24<=w_1_472; wr25<=w_1_473; wr26<=w_1_474; wr27<=w_1_475; wr28<=w_1_476; wr29<=w_1_477; wr30<=w_1_478; wr31<=w_1_479; wr32<=w_1_480; wr33<=w_1_481; wr34<=w_1_482; wr35<=w_1_483; wr36<=w_1_484; wr37<=w_1_485; wr38<=w_1_486; wr39<=w_1_487; wr40<=w_1_488; wr41<=w_1_489; wr42<=w_1_490; wr43<=w_1_491; wr44<=w_1_492; wr45<=w_1_493; wr46<=w_1_494; wr47<=w_1_495; wr48<=w_1_496; wr49<=w_1_497; wr50<=w_1_498; wr51<=w_1_499; wr52<=w_1_500; wr53<=w_1_501; wr54<=w_1_502; wr55<=w_1_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd25:
					begin
						wr0<=w_1_504; wr1<=w_1_505; wr2<=w_1_506; wr3<=w_1_507; wr4<=w_1_508; wr5<=w_1_509; wr6<=w_1_510; wr7<=w_1_511; wr8<=w_1_512; wr9<=w_1_513; wr10<=w_1_514; wr11<=w_1_515; wr12<=w_1_516; wr13<=w_1_517; wr14<=w_1_518; wr15<=w_1_519; wr16<=w_1_520; wr17<=w_1_521; wr18<=w_1_522; wr19<=w_1_523; wr20<=w_1_524; wr21<=w_1_525; wr22<=w_1_526; wr23<=w_1_527; wr24<=w_1_528; wr25<=w_1_529; wr26<=w_1_530; wr27<=w_1_531; wr28<=w_1_532; wr29<=w_1_533; wr30<=w_1_534; wr31<=w_1_535; wr32<=w_1_536; wr33<=w_1_537; wr34<=w_1_538; wr35<=w_1_539; wr36<=w_1_540; wr37<=w_1_541; wr38<=w_1_542; wr39<=w_1_543; wr40<=w_1_544; wr41<=w_1_545; wr42<=w_1_546; wr43<=w_1_547; wr44<=w_1_548; wr45<=w_1_549; wr46<=w_1_550; wr47<=w_1_551; wr48<=w_1_552; wr49<=w_1_553; wr50<=w_1_554; wr51<=w_1_555; wr52<=w_1_556; wr53<=w_1_557; wr54<=w_1_558; wr55<=w_1_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd26:
					begin
						wr0<=w_1_560; wr1<=w_1_561; wr2<=w_1_562; wr3<=w_1_563; wr4<=w_1_564; wr5<=w_1_565; wr6<=w_1_566; wr7<=w_1_567; wr8<=w_1_568; wr9<=w_1_569; wr10<=w_1_570; wr11<=w_1_571; wr12<=w_1_572; wr13<=w_1_573; wr14<=w_1_574; wr15<=w_1_575; wr16<=w_1_576; wr17<=w_1_577; wr18<=w_1_578; wr19<=w_1_579; wr20<=w_1_580; wr21<=w_1_581; wr22<=w_1_582; wr23<=w_1_583; wr24<=w_1_584; wr25<=w_1_585; wr26<=w_1_586; wr27<=w_1_587; wr28<=w_1_588; wr29<=w_1_589; wr30<=w_1_590; wr31<=w_1_591; wr32<=w_1_592; wr33<=w_1_593; wr34<=w_1_594; wr35<=w_1_595; wr36<=w_1_596; wr37<=w_1_597; wr38<=w_1_598; wr39<=w_1_599; wr40<=w_1_600; wr41<=w_1_601; wr42<=w_1_602; wr43<=w_1_603; wr44<=w_1_604; wr45<=w_1_605; wr46<=w_1_606; wr47<=w_1_607; wr48<=w_1_608; wr49<=w_1_609; wr50<=w_1_610; wr51<=w_1_611; wr52<=w_1_612; wr53<=w_1_613; wr54<=w_1_614; wr55<=w_1_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd27:
					begin
						wr0<=w_1_616; wr1<=w_1_617; wr2<=w_1_618; wr3<=w_1_619; wr4<=w_1_620; wr5<=w_1_621; wr6<=w_1_622; wr7<=w_1_623; wr8<=w_1_624; wr9<=w_1_625; wr10<=w_1_626; wr11<=w_1_627; wr12<=w_1_628; wr13<=w_1_629; wr14<=w_1_630; wr15<=w_1_631; wr16<=w_1_632; wr17<=w_1_633; wr18<=w_1_634; wr19<=w_1_635; wr20<=w_1_636; wr21<=w_1_637; wr22<=w_1_638; wr23<=w_1_639; wr24<=w_1_640; wr25<=w_1_641; wr26<=w_1_642; wr27<=w_1_643; wr28<=w_1_644; wr29<=w_1_645; wr30<=w_1_646; wr31<=w_1_647; wr32<=w_1_648; wr33<=w_1_649; wr34<=w_1_650; wr35<=w_1_651; wr36<=w_1_652; wr37<=w_1_653; wr38<=w_1_654; wr39<=w_1_655; wr40<=w_1_656; wr41<=w_1_657; wr42<=w_1_658; wr43<=w_1_659; wr44<=w_1_660; wr45<=w_1_661; wr46<=w_1_662; wr47<=w_1_663; wr48<=w_1_664; wr49<=w_1_665; wr50<=w_1_666; wr51<=w_1_667; wr52<=w_1_668; wr53<=w_1_669; wr54<=w_1_670; wr55<=w_1_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd28:
					begin
						wr0<=w_1_672; wr1<=w_1_673; wr2<=w_1_674; wr3<=w_1_675; wr4<=w_1_676; wr5<=w_1_677; wr6<=w_1_678; wr7<=w_1_679; wr8<=w_1_680; wr9<=w_1_681; wr10<=w_1_682; wr11<=w_1_683; wr12<=w_1_684; wr13<=w_1_685; wr14<=w_1_686; wr15<=w_1_687; wr16<=w_1_688; wr17<=w_1_689; wr18<=w_1_690; wr19<=w_1_691; wr20<=w_1_692; wr21<=w_1_693; wr22<=w_1_694; wr23<=w_1_695; wr24<=w_1_696; wr25<=w_1_697; wr26<=w_1_698; wr27<=w_1_699; wr28<=w_1_700; wr29<=w_1_701; wr30<=w_1_702; wr31<=w_1_703; wr32<=w_1_704; wr33<=w_1_705; wr34<=w_1_706; wr35<=w_1_707; wr36<=w_1_708; wr37<=w_1_709; wr38<=w_1_710; wr39<=w_1_711; wr40<=w_1_712; wr41<=w_1_713; wr42<=w_1_714; wr43<=w_1_715; wr44<=w_1_716; wr45<=w_1_717; wr46<=w_1_718; wr47<=w_1_719; wr48<=w_1_720; wr49<=w_1_721; wr50<=w_1_722; wr51<=w_1_723; wr52<=w_1_724; wr53<=w_1_725; wr54<=w_1_726; wr55<=w_1_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd29:
					begin
						wr0<=w_1_728; wr1<=w_1_729; wr2<=w_1_730; wr3<=w_1_731; wr4<=w_1_732; wr5<=w_1_733; wr6<=w_1_734; wr7<=w_1_735; wr8<=w_1_736; wr9<=w_1_737; wr10<=w_1_738; wr11<=w_1_739; wr12<=w_1_740; wr13<=w_1_741; wr14<=w_1_742; wr15<=w_1_743; wr16<=w_1_744; wr17<=w_1_745; wr18<=w_1_746; wr19<=w_1_747; wr20<=w_1_748; wr21<=w_1_749; wr22<=w_1_750; wr23<=w_1_751; wr24<=w_1_752; wr25<=w_1_753; wr26<=w_1_754; wr27<=w_1_755; wr28<=w_1_756; wr29<=w_1_757; wr30<=w_1_758; wr31<=w_1_759; wr32<=w_1_760; wr33<=w_1_761; wr34<=w_1_762; wr35<=w_1_763; wr36<=w_1_764; wr37<=w_1_765; wr38<=w_1_766; wr39<=w_1_767; wr40<=w_1_768; wr41<=w_1_769; wr42<=w_1_770; wr43<=w_1_771; wr44<=w_1_772; wr45<=w_1_773; wr46<=w_1_774; wr47<=w_1_775; wr48<=w_1_776; wr49<=w_1_777; wr50<=w_1_778; wr51<=w_1_779; wr52<=w_1_780; wr53<=w_1_781; wr54<=w_1_782; wr55<=w_1_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd30:
					begin
						bias_p<=px_784;
						bias_w<=w_1_784;
						select<=select+1;
					end
				8'd31:
					begin
						wr0<=w_2_0; wr1<=w_2_1; wr2<=w_2_2; wr3<=w_2_3; wr4<=w_2_4; wr5<=w_2_5; wr6<=w_2_6; wr7<=w_2_7; wr8<=w_2_8; wr9<=w_2_9; wr10<=w_2_10; wr11<=w_2_11; wr12<=w_2_12; wr13<=w_2_13; wr14<=w_2_14; wr15<=w_2_15; wr16<=w_2_16; wr17<=w_2_17; wr18<=w_2_18; wr19<=w_2_19; wr20<=w_2_20; wr21<=w_2_21; wr22<=w_2_22; wr23<=w_2_23; wr24<=w_2_24; wr25<=w_2_25; wr26<=w_2_26; wr27<=w_2_27; wr28<=w_2_28; wr29<=w_2_29; wr30<=w_2_30; wr31<=w_2_31; wr32<=w_2_32; wr33<=w_2_33; wr34<=w_2_34; wr35<=w_2_35; wr36<=w_2_36; wr37<=w_2_37; wr38<=w_2_38; wr39<=w_2_39; wr40<=w_2_40; wr41<=w_2_41; wr42<=w_2_42; wr43<=w_2_43; wr44<=w_2_44; wr45<=w_2_45; wr46<=w_2_46; wr47<=w_2_47; wr48<=w_2_48; wr49<=w_2_49; wr50<=w_2_50; wr51<=w_2_51; wr52<=w_2_52; wr53<=w_2_53; wr54<=w_2_54; wr55<=w_2_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd32:
					begin
						wr0<=w_2_56; wr1<=w_2_57; wr2<=w_2_58; wr3<=w_2_59; wr4<=w_2_60; wr5<=w_2_61; wr6<=w_2_62; wr7<=w_2_63; wr8<=w_2_64; wr9<=w_2_65; wr10<=w_2_66; wr11<=w_2_67; wr12<=w_2_68; wr13<=w_2_69; wr14<=w_2_70; wr15<=w_2_71; wr16<=w_2_72; wr17<=w_2_73; wr18<=w_2_74; wr19<=w_2_75; wr20<=w_2_76; wr21<=w_2_77; wr22<=w_2_78; wr23<=w_2_79; wr24<=w_2_80; wr25<=w_2_81; wr26<=w_2_82; wr27<=w_2_83; wr28<=w_2_84; wr29<=w_2_85; wr30<=w_2_86; wr31<=w_2_87; wr32<=w_2_88; wr33<=w_2_89; wr34<=w_2_90; wr35<=w_2_91; wr36<=w_2_92; wr37<=w_2_93; wr38<=w_2_94; wr39<=w_2_95; wr40<=w_2_96; wr41<=w_2_97; wr42<=w_2_98; wr43<=w_2_99; wr44<=w_2_100; wr45<=w_2_101; wr46<=w_2_102; wr47<=w_2_103; wr48<=w_2_104; wr49<=w_2_105; wr50<=w_2_106; wr51<=w_2_107; wr52<=w_2_108; wr53<=w_2_109; wr54<=w_2_110; wr55<=w_2_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd33:
					begin
						wr0<=w_2_112; wr1<=w_2_113; wr2<=w_2_114; wr3<=w_2_115; wr4<=w_2_116; wr5<=w_2_117; wr6<=w_2_118; wr7<=w_2_119; wr8<=w_2_120; wr9<=w_2_121; wr10<=w_2_122; wr11<=w_2_123; wr12<=w_2_124; wr13<=w_2_125; wr14<=w_2_126; wr15<=w_2_127; wr16<=w_2_128; wr17<=w_2_129; wr18<=w_2_130; wr19<=w_2_131; wr20<=w_2_132; wr21<=w_2_133; wr22<=w_2_134; wr23<=w_2_135; wr24<=w_2_136; wr25<=w_2_137; wr26<=w_2_138; wr27<=w_2_139; wr28<=w_2_140; wr29<=w_2_141; wr30<=w_2_142; wr31<=w_2_143; wr32<=w_2_144; wr33<=w_2_145; wr34<=w_2_146; wr35<=w_2_147; wr36<=w_2_148; wr37<=w_2_149; wr38<=w_2_150; wr39<=w_2_151; wr40<=w_2_152; wr41<=w_2_153; wr42<=w_2_154; wr43<=w_2_155; wr44<=w_2_156; wr45<=w_2_157; wr46<=w_2_158; wr47<=w_2_159; wr48<=w_2_160; wr49<=w_2_161; wr50<=w_2_162; wr51<=w_2_163; wr52<=w_2_164; wr53<=w_2_165; wr54<=w_2_166; wr55<=w_2_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd34:
					begin
						wr0<=w_2_168; wr1<=w_2_169; wr2<=w_2_170; wr3<=w_2_171; wr4<=w_2_172; wr5<=w_2_173; wr6<=w_2_174; wr7<=w_2_175; wr8<=w_2_176; wr9<=w_2_177; wr10<=w_2_178; wr11<=w_2_179; wr12<=w_2_180; wr13<=w_2_181; wr14<=w_2_182; wr15<=w_2_183; wr16<=w_2_184; wr17<=w_2_185; wr18<=w_2_186; wr19<=w_2_187; wr20<=w_2_188; wr21<=w_2_189; wr22<=w_2_190; wr23<=w_2_191; wr24<=w_2_192; wr25<=w_2_193; wr26<=w_2_194; wr27<=w_2_195; wr28<=w_2_196; wr29<=w_2_197; wr30<=w_2_198; wr31<=w_2_199; wr32<=w_2_200; wr33<=w_2_201; wr34<=w_2_202; wr35<=w_2_203; wr36<=w_2_204; wr37<=w_2_205; wr38<=w_2_206; wr39<=w_2_207; wr40<=w_2_208; wr41<=w_2_209; wr42<=w_2_210; wr43<=w_2_211; wr44<=w_2_212; wr45<=w_2_213; wr46<=w_2_214; wr47<=w_2_215; wr48<=w_2_216; wr49<=w_2_217; wr50<=w_2_218; wr51<=w_2_219; wr52<=w_2_220; wr53<=w_2_221; wr54<=w_2_222; wr55<=w_2_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd35:
					begin
						wr0<=w_2_224; wr1<=w_2_225; wr2<=w_2_226; wr3<=w_2_227; wr4<=w_2_228; wr5<=w_2_229; wr6<=w_2_230; wr7<=w_2_231; wr8<=w_2_232; wr9<=w_2_233; wr10<=w_2_234; wr11<=w_2_235; wr12<=w_2_236; wr13<=w_2_237; wr14<=w_2_238; wr15<=w_2_239; wr16<=w_2_240; wr17<=w_2_241; wr18<=w_2_242; wr19<=w_2_243; wr20<=w_2_244; wr21<=w_2_245; wr22<=w_2_246; wr23<=w_2_247; wr24<=w_2_248; wr25<=w_2_249; wr26<=w_2_250; wr27<=w_2_251; wr28<=w_2_252; wr29<=w_2_253; wr30<=w_2_254; wr31<=w_2_255; wr32<=w_2_256; wr33<=w_2_257; wr34<=w_2_258; wr35<=w_2_259; wr36<=w_2_260; wr37<=w_2_261; wr38<=w_2_262; wr39<=w_2_263; wr40<=w_2_264; wr41<=w_2_265; wr42<=w_2_266; wr43<=w_2_267; wr44<=w_2_268; wr45<=w_2_269; wr46<=w_2_270; wr47<=w_2_271; wr48<=w_2_272; wr49<=w_2_273; wr50<=w_2_274; wr51<=w_2_275; wr52<=w_2_276; wr53<=w_2_277; wr54<=w_2_278; wr55<=w_2_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd36:
					begin
						wr0<=w_2_280; wr1<=w_2_281; wr2<=w_2_282; wr3<=w_2_283; wr4<=w_2_284; wr5<=w_2_285; wr6<=w_2_286; wr7<=w_2_287; wr8<=w_2_288; wr9<=w_2_289; wr10<=w_2_290; wr11<=w_2_291; wr12<=w_2_292; wr13<=w_2_293; wr14<=w_2_294; wr15<=w_2_295; wr16<=w_2_296; wr17<=w_2_297; wr18<=w_2_298; wr19<=w_2_299; wr20<=w_2_300; wr21<=w_2_301; wr22<=w_2_302; wr23<=w_2_303; wr24<=w_2_304; wr25<=w_2_305; wr26<=w_2_306; wr27<=w_2_307; wr28<=w_2_308; wr29<=w_2_309; wr30<=w_2_310; wr31<=w_2_311; wr32<=w_2_312; wr33<=w_2_313; wr34<=w_2_314; wr35<=w_2_315; wr36<=w_2_316; wr37<=w_2_317; wr38<=w_2_318; wr39<=w_2_319; wr40<=w_2_320; wr41<=w_2_321; wr42<=w_2_322; wr43<=w_2_323; wr44<=w_2_324; wr45<=w_2_325; wr46<=w_2_326; wr47<=w_2_327; wr48<=w_2_328; wr49<=w_2_329; wr50<=w_2_330; wr51<=w_2_331; wr52<=w_2_332; wr53<=w_2_333; wr54<=w_2_334; wr55<=w_2_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd37:
					begin
						wr0<=w_2_336; wr1<=w_2_337; wr2<=w_2_338; wr3<=w_2_339; wr4<=w_2_340; wr5<=w_2_341; wr6<=w_2_342; wr7<=w_2_343; wr8<=w_2_344; wr9<=w_2_345; wr10<=w_2_346; wr11<=w_2_347; wr12<=w_2_348; wr13<=w_2_349; wr14<=w_2_350; wr15<=w_2_351; wr16<=w_2_352; wr17<=w_2_353; wr18<=w_2_354; wr19<=w_2_355; wr20<=w_2_356; wr21<=w_2_357; wr22<=w_2_358; wr23<=w_2_359; wr24<=w_2_360; wr25<=w_2_361; wr26<=w_2_362; wr27<=w_2_363; wr28<=w_2_364; wr29<=w_2_365; wr30<=w_2_366; wr31<=w_2_367; wr32<=w_2_368; wr33<=w_2_369; wr34<=w_2_370; wr35<=w_2_371; wr36<=w_2_372; wr37<=w_2_373; wr38<=w_2_374; wr39<=w_2_375; wr40<=w_2_376; wr41<=w_2_377; wr42<=w_2_378; wr43<=w_2_379; wr44<=w_2_380; wr45<=w_2_381; wr46<=w_2_382; wr47<=w_2_383; wr48<=w_2_384; wr49<=w_2_385; wr50<=w_2_386; wr51<=w_2_387; wr52<=w_2_388; wr53<=w_2_389; wr54<=w_2_390; wr55<=w_2_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd38:
					begin
						wr0<=w_2_392; wr1<=w_2_393; wr2<=w_2_394; wr3<=w_2_395; wr4<=w_2_396; wr5<=w_2_397; wr6<=w_2_398; wr7<=w_2_399; wr8<=w_2_400; wr9<=w_2_401; wr10<=w_2_402; wr11<=w_2_403; wr12<=w_2_404; wr13<=w_2_405; wr14<=w_2_406; wr15<=w_2_407; wr16<=w_2_408; wr17<=w_2_409; wr18<=w_2_410; wr19<=w_2_411; wr20<=w_2_412; wr21<=w_2_413; wr22<=w_2_414; wr23<=w_2_415; wr24<=w_2_416; wr25<=w_2_417; wr26<=w_2_418; wr27<=w_2_419; wr28<=w_2_420; wr29<=w_2_421; wr30<=w_2_422; wr31<=w_2_423; wr32<=w_2_424; wr33<=w_2_425; wr34<=w_2_426; wr35<=w_2_427; wr36<=w_2_428; wr37<=w_2_429; wr38<=w_2_430; wr39<=w_2_431; wr40<=w_2_432; wr41<=w_2_433; wr42<=w_2_434; wr43<=w_2_435; wr44<=w_2_436; wr45<=w_2_437; wr46<=w_2_438; wr47<=w_2_439; wr48<=w_2_440; wr49<=w_2_441; wr50<=w_2_442; wr51<=w_2_443; wr52<=w_2_444; wr53<=w_2_445; wr54<=w_2_446; wr55<=w_2_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd39:
					begin
						wr0<=w_2_448; wr1<=w_2_449; wr2<=w_2_450; wr3<=w_2_451; wr4<=w_2_452; wr5<=w_2_453; wr6<=w_2_454; wr7<=w_2_455; wr8<=w_2_456; wr9<=w_2_457; wr10<=w_2_458; wr11<=w_2_459; wr12<=w_2_460; wr13<=w_2_461; wr14<=w_2_462; wr15<=w_2_463; wr16<=w_2_464; wr17<=w_2_465; wr18<=w_2_466; wr19<=w_2_467; wr20<=w_2_468; wr21<=w_2_469; wr22<=w_2_470; wr23<=w_2_471; wr24<=w_2_472; wr25<=w_2_473; wr26<=w_2_474; wr27<=w_2_475; wr28<=w_2_476; wr29<=w_2_477; wr30<=w_2_478; wr31<=w_2_479; wr32<=w_2_480; wr33<=w_2_481; wr34<=w_2_482; wr35<=w_2_483; wr36<=w_2_484; wr37<=w_2_485; wr38<=w_2_486; wr39<=w_2_487; wr40<=w_2_488; wr41<=w_2_489; wr42<=w_2_490; wr43<=w_2_491; wr44<=w_2_492; wr45<=w_2_493; wr46<=w_2_494; wr47<=w_2_495; wr48<=w_2_496; wr49<=w_2_497; wr50<=w_2_498; wr51<=w_2_499; wr52<=w_2_500; wr53<=w_2_501; wr54<=w_2_502; wr55<=w_2_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd40:
					begin
						wr0<=w_2_504; wr1<=w_2_505; wr2<=w_2_506; wr3<=w_2_507; wr4<=w_2_508; wr5<=w_2_509; wr6<=w_2_510; wr7<=w_2_511; wr8<=w_2_512; wr9<=w_2_513; wr10<=w_2_514; wr11<=w_2_515; wr12<=w_2_516; wr13<=w_2_517; wr14<=w_2_518; wr15<=w_2_519; wr16<=w_2_520; wr17<=w_2_521; wr18<=w_2_522; wr19<=w_2_523; wr20<=w_2_524; wr21<=w_2_525; wr22<=w_2_526; wr23<=w_2_527; wr24<=w_2_528; wr25<=w_2_529; wr26<=w_2_530; wr27<=w_2_531; wr28<=w_2_532; wr29<=w_2_533; wr30<=w_2_534; wr31<=w_2_535; wr32<=w_2_536; wr33<=w_2_537; wr34<=w_2_538; wr35<=w_2_539; wr36<=w_2_540; wr37<=w_2_541; wr38<=w_2_542; wr39<=w_2_543; wr40<=w_2_544; wr41<=w_2_545; wr42<=w_2_546; wr43<=w_2_547; wr44<=w_2_548; wr45<=w_2_549; wr46<=w_2_550; wr47<=w_2_551; wr48<=w_2_552; wr49<=w_2_553; wr50<=w_2_554; wr51<=w_2_555; wr52<=w_2_556; wr53<=w_2_557; wr54<=w_2_558; wr55<=w_2_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd41:
					begin
						wr0<=w_2_560; wr1<=w_2_561; wr2<=w_2_562; wr3<=w_2_563; wr4<=w_2_564; wr5<=w_2_565; wr6<=w_2_566; wr7<=w_2_567; wr8<=w_2_568; wr9<=w_2_569; wr10<=w_2_570; wr11<=w_2_571; wr12<=w_2_572; wr13<=w_2_573; wr14<=w_2_574; wr15<=w_2_575; wr16<=w_2_576; wr17<=w_2_577; wr18<=w_2_578; wr19<=w_2_579; wr20<=w_2_580; wr21<=w_2_581; wr22<=w_2_582; wr23<=w_2_583; wr24<=w_2_584; wr25<=w_2_585; wr26<=w_2_586; wr27<=w_2_587; wr28<=w_2_588; wr29<=w_2_589; wr30<=w_2_590; wr31<=w_2_591; wr32<=w_2_592; wr33<=w_2_593; wr34<=w_2_594; wr35<=w_2_595; wr36<=w_2_596; wr37<=w_2_597; wr38<=w_2_598; wr39<=w_2_599; wr40<=w_2_600; wr41<=w_2_601; wr42<=w_2_602; wr43<=w_2_603; wr44<=w_2_604; wr45<=w_2_605; wr46<=w_2_606; wr47<=w_2_607; wr48<=w_2_608; wr49<=w_2_609; wr50<=w_2_610; wr51<=w_2_611; wr52<=w_2_612; wr53<=w_2_613; wr54<=w_2_614; wr55<=w_2_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd42:
					begin
						wr0<=w_2_616; wr1<=w_2_617; wr2<=w_2_618; wr3<=w_2_619; wr4<=w_2_620; wr5<=w_2_621; wr6<=w_2_622; wr7<=w_2_623; wr8<=w_2_624; wr9<=w_2_625; wr10<=w_2_626; wr11<=w_2_627; wr12<=w_2_628; wr13<=w_2_629; wr14<=w_2_630; wr15<=w_2_631; wr16<=w_2_632; wr17<=w_2_633; wr18<=w_2_634; wr19<=w_2_635; wr20<=w_2_636; wr21<=w_2_637; wr22<=w_2_638; wr23<=w_2_639; wr24<=w_2_640; wr25<=w_2_641; wr26<=w_2_642; wr27<=w_2_643; wr28<=w_2_644; wr29<=w_2_645; wr30<=w_2_646; wr31<=w_2_647; wr32<=w_2_648; wr33<=w_2_649; wr34<=w_2_650; wr35<=w_2_651; wr36<=w_2_652; wr37<=w_2_653; wr38<=w_2_654; wr39<=w_2_655; wr40<=w_2_656; wr41<=w_2_657; wr42<=w_2_658; wr43<=w_2_659; wr44<=w_2_660; wr45<=w_2_661; wr46<=w_2_662; wr47<=w_2_663; wr48<=w_2_664; wr49<=w_2_665; wr50<=w_2_666; wr51<=w_2_667; wr52<=w_2_668; wr53<=w_2_669; wr54<=w_2_670; wr55<=w_2_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd43:
					begin
						wr0<=w_2_672; wr1<=w_2_673; wr2<=w_2_674; wr3<=w_2_675; wr4<=w_2_676; wr5<=w_2_677; wr6<=w_2_678; wr7<=w_2_679; wr8<=w_2_680; wr9<=w_2_681; wr10<=w_2_682; wr11<=w_2_683; wr12<=w_2_684; wr13<=w_2_685; wr14<=w_2_686; wr15<=w_2_687; wr16<=w_2_688; wr17<=w_2_689; wr18<=w_2_690; wr19<=w_2_691; wr20<=w_2_692; wr21<=w_2_693; wr22<=w_2_694; wr23<=w_2_695; wr24<=w_2_696; wr25<=w_2_697; wr26<=w_2_698; wr27<=w_2_699; wr28<=w_2_700; wr29<=w_2_701; wr30<=w_2_702; wr31<=w_2_703; wr32<=w_2_704; wr33<=w_2_705; wr34<=w_2_706; wr35<=w_2_707; wr36<=w_2_708; wr37<=w_2_709; wr38<=w_2_710; wr39<=w_2_711; wr40<=w_2_712; wr41<=w_2_713; wr42<=w_2_714; wr43<=w_2_715; wr44<=w_2_716; wr45<=w_2_717; wr46<=w_2_718; wr47<=w_2_719; wr48<=w_2_720; wr49<=w_2_721; wr50<=w_2_722; wr51<=w_2_723; wr52<=w_2_724; wr53<=w_2_725; wr54<=w_2_726; wr55<=w_2_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd44:
					begin
						wr0<=w_2_728; wr1<=w_2_729; wr2<=w_2_730; wr3<=w_2_731; wr4<=w_2_732; wr5<=w_2_733; wr6<=w_2_734; wr7<=w_2_735; wr8<=w_2_736; wr9<=w_2_737; wr10<=w_2_738; wr11<=w_2_739; wr12<=w_2_740; wr13<=w_2_741; wr14<=w_2_742; wr15<=w_2_743; wr16<=w_2_744; wr17<=w_2_745; wr18<=w_2_746; wr19<=w_2_747; wr20<=w_2_748; wr21<=w_2_749; wr22<=w_2_750; wr23<=w_2_751; wr24<=w_2_752; wr25<=w_2_753; wr26<=w_2_754; wr27<=w_2_755; wr28<=w_2_756; wr29<=w_2_757; wr30<=w_2_758; wr31<=w_2_759; wr32<=w_2_760; wr33<=w_2_761; wr34<=w_2_762; wr35<=w_2_763; wr36<=w_2_764; wr37<=w_2_765; wr38<=w_2_766; wr39<=w_2_767; wr40<=w_2_768; wr41<=w_2_769; wr42<=w_2_770; wr43<=w_2_771; wr44<=w_2_772; wr45<=w_2_773; wr46<=w_2_774; wr47<=w_2_775; wr48<=w_2_776; wr49<=w_2_777; wr50<=w_2_778; wr51<=w_2_779; wr52<=w_2_780; wr53<=w_2_781; wr54<=w_2_782; wr55<=w_2_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd45:
					begin
						bias_p<=px_784;
						bias_w<=w_2_784;
						select<=select+1;
						
					end
				8'd46:
					begin
						wr0<=w_3_0; wr1<=w_3_1; wr2<=w_3_2; wr3<=w_3_3; wr4<=w_3_4; wr5<=w_3_5; wr6<=w_3_6; wr7<=w_3_7; wr8<=w_3_8; wr9<=w_3_9; wr10<=w_3_10; wr11<=w_3_11; wr12<=w_3_12; wr13<=w_3_13; wr14<=w_3_14; wr15<=w_3_15; wr16<=w_3_16; wr17<=w_3_17; wr18<=w_3_18; wr19<=w_3_19; wr20<=w_3_20; wr21<=w_3_21; wr22<=w_3_22; wr23<=w_3_23; wr24<=w_3_24; wr25<=w_3_25; wr26<=w_3_26; wr27<=w_3_27; wr28<=w_3_28; wr29<=w_3_29; wr30<=w_3_30; wr31<=w_3_31; wr32<=w_3_32; wr33<=w_3_33; wr34<=w_3_34; wr35<=w_3_35; wr36<=w_3_36; wr37<=w_3_37; wr38<=w_3_38; wr39<=w_3_39; wr40<=w_3_40; wr41<=w_3_41; wr42<=w_3_42; wr43<=w_3_43; wr44<=w_3_44; wr45<=w_3_45; wr46<=w_3_46; wr47<=w_3_47; wr48<=w_3_48; wr49<=w_3_49; wr50<=w_3_50; wr51<=w_3_51; wr52<=w_3_52; wr53<=w_3_53; wr54<=w_3_54; wr55<=w_3_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd47:
					begin
						wr0<=w_3_56; wr1<=w_3_57; wr2<=w_3_58; wr3<=w_3_59; wr4<=w_3_60; wr5<=w_3_61; wr6<=w_3_62; wr7<=w_3_63; wr8<=w_3_64; wr9<=w_3_65; wr10<=w_3_66; wr11<=w_3_67; wr12<=w_3_68; wr13<=w_3_69; wr14<=w_3_70; wr15<=w_3_71; wr16<=w_3_72; wr17<=w_3_73; wr18<=w_3_74; wr19<=w_3_75; wr20<=w_3_76; wr21<=w_3_77; wr22<=w_3_78; wr23<=w_3_79; wr24<=w_3_80; wr25<=w_3_81; wr26<=w_3_82; wr27<=w_3_83; wr28<=w_3_84; wr29<=w_3_85; wr30<=w_3_86; wr31<=w_3_87; wr32<=w_3_88; wr33<=w_3_89; wr34<=w_3_90; wr35<=w_3_91; wr36<=w_3_92; wr37<=w_3_93; wr38<=w_3_94; wr39<=w_3_95; wr40<=w_3_96; wr41<=w_3_97; wr42<=w_3_98; wr43<=w_3_99; wr44<=w_3_100; wr45<=w_3_101; wr46<=w_3_102; wr47<=w_3_103; wr48<=w_3_104; wr49<=w_3_105; wr50<=w_3_106; wr51<=w_3_107; wr52<=w_3_108; wr53<=w_3_109; wr54<=w_3_110; wr55<=w_3_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd48:
					begin
						wr0<=w_3_112; wr1<=w_3_113; wr2<=w_3_114; wr3<=w_3_115; wr4<=w_3_116; wr5<=w_3_117; wr6<=w_3_118; wr7<=w_3_119; wr8<=w_3_120; wr9<=w_3_121; wr10<=w_3_122; wr11<=w_3_123; wr12<=w_3_124; wr13<=w_3_125; wr14<=w_3_126; wr15<=w_3_127; wr16<=w_3_128; wr17<=w_3_129; wr18<=w_3_130; wr19<=w_3_131; wr20<=w_3_132; wr21<=w_3_133; wr22<=w_3_134; wr23<=w_3_135; wr24<=w_3_136; wr25<=w_3_137; wr26<=w_3_138; wr27<=w_3_139; wr28<=w_3_140; wr29<=w_3_141; wr30<=w_3_142; wr31<=w_3_143; wr32<=w_3_144; wr33<=w_3_145; wr34<=w_3_146; wr35<=w_3_147; wr36<=w_3_148; wr37<=w_3_149; wr38<=w_3_150; wr39<=w_3_151; wr40<=w_3_152; wr41<=w_3_153; wr42<=w_3_154; wr43<=w_3_155; wr44<=w_3_156; wr45<=w_3_157; wr46<=w_3_158; wr47<=w_3_159; wr48<=w_3_160; wr49<=w_3_161; wr50<=w_3_162; wr51<=w_3_163; wr52<=w_3_164; wr53<=w_3_165; wr54<=w_3_166; wr55<=w_3_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd49:
					begin
						wr0<=w_3_168; wr1<=w_3_169; wr2<=w_3_170; wr3<=w_3_171; wr4<=w_3_172; wr5<=w_3_173; wr6<=w_3_174; wr7<=w_3_175; wr8<=w_3_176; wr9<=w_3_177; wr10<=w_3_178; wr11<=w_3_179; wr12<=w_3_180; wr13<=w_3_181; wr14<=w_3_182; wr15<=w_3_183; wr16<=w_3_184; wr17<=w_3_185; wr18<=w_3_186; wr19<=w_3_187; wr20<=w_3_188; wr21<=w_3_189; wr22<=w_3_190; wr23<=w_3_191; wr24<=w_3_192; wr25<=w_3_193; wr26<=w_3_194; wr27<=w_3_195; wr28<=w_3_196; wr29<=w_3_197; wr30<=w_3_198; wr31<=w_3_199; wr32<=w_3_200; wr33<=w_3_201; wr34<=w_3_202; wr35<=w_3_203; wr36<=w_3_204; wr37<=w_3_205; wr38<=w_3_206; wr39<=w_3_207; wr40<=w_3_208; wr41<=w_3_209; wr42<=w_3_210; wr43<=w_3_211; wr44<=w_3_212; wr45<=w_3_213; wr46<=w_3_214; wr47<=w_3_215; wr48<=w_3_216; wr49<=w_3_217; wr50<=w_3_218; wr51<=w_3_219; wr52<=w_3_220; wr53<=w_3_221; wr54<=w_3_222; wr55<=w_3_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd50:
					begin
						wr0<=w_3_224; wr1<=w_3_225; wr2<=w_3_226; wr3<=w_3_227; wr4<=w_3_228; wr5<=w_3_229; wr6<=w_3_230; wr7<=w_3_231; wr8<=w_3_232; wr9<=w_3_233; wr10<=w_3_234; wr11<=w_3_235; wr12<=w_3_236; wr13<=w_3_237; wr14<=w_3_238; wr15<=w_3_239; wr16<=w_3_240; wr17<=w_3_241; wr18<=w_3_242; wr19<=w_3_243; wr20<=w_3_244; wr21<=w_3_245; wr22<=w_3_246; wr23<=w_3_247; wr24<=w_3_248; wr25<=w_3_249; wr26<=w_3_250; wr27<=w_3_251; wr28<=w_3_252; wr29<=w_3_253; wr30<=w_3_254; wr31<=w_3_255; wr32<=w_3_256; wr33<=w_3_257; wr34<=w_3_258; wr35<=w_3_259; wr36<=w_3_260; wr37<=w_3_261; wr38<=w_3_262; wr39<=w_3_263; wr40<=w_3_264; wr41<=w_3_265; wr42<=w_3_266; wr43<=w_3_267; wr44<=w_3_268; wr45<=w_3_269; wr46<=w_3_270; wr47<=w_3_271; wr48<=w_3_272; wr49<=w_3_273; wr50<=w_3_274; wr51<=w_3_275; wr52<=w_3_276; wr53<=w_3_277; wr54<=w_3_278; wr55<=w_3_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd51:
					begin
						wr0<=w_3_280; wr1<=w_3_281; wr2<=w_3_282; wr3<=w_3_283; wr4<=w_3_284; wr5<=w_3_285; wr6<=w_3_286; wr7<=w_3_287; wr8<=w_3_288; wr9<=w_3_289; wr10<=w_3_290; wr11<=w_3_291; wr12<=w_3_292; wr13<=w_3_293; wr14<=w_3_294; wr15<=w_3_295; wr16<=w_3_296; wr17<=w_3_297; wr18<=w_3_298; wr19<=w_3_299; wr20<=w_3_300; wr21<=w_3_301; wr22<=w_3_302; wr23<=w_3_303; wr24<=w_3_304; wr25<=w_3_305; wr26<=w_3_306; wr27<=w_3_307; wr28<=w_3_308; wr29<=w_3_309; wr30<=w_3_310; wr31<=w_3_311; wr32<=w_3_312; wr33<=w_3_313; wr34<=w_3_314; wr35<=w_3_315; wr36<=w_3_316; wr37<=w_3_317; wr38<=w_3_318; wr39<=w_3_319; wr40<=w_3_320; wr41<=w_3_321; wr42<=w_3_322; wr43<=w_3_323; wr44<=w_3_324; wr45<=w_3_325; wr46<=w_3_326; wr47<=w_3_327; wr48<=w_3_328; wr49<=w_3_329; wr50<=w_3_330; wr51<=w_3_331; wr52<=w_3_332; wr53<=w_3_333; wr54<=w_3_334; wr55<=w_3_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd52:
					begin
						wr0<=w_3_336; wr1<=w_3_337; wr2<=w_3_338; wr3<=w_3_339; wr4<=w_3_340; wr5<=w_3_341; wr6<=w_3_342; wr7<=w_3_343; wr8<=w_3_344; wr9<=w_3_345; wr10<=w_3_346; wr11<=w_3_347; wr12<=w_3_348; wr13<=w_3_349; wr14<=w_3_350; wr15<=w_3_351; wr16<=w_3_352; wr17<=w_3_353; wr18<=w_3_354; wr19<=w_3_355; wr20<=w_3_356; wr21<=w_3_357; wr22<=w_3_358; wr23<=w_3_359; wr24<=w_3_360; wr25<=w_3_361; wr26<=w_3_362; wr27<=w_3_363; wr28<=w_3_364; wr29<=w_3_365; wr30<=w_3_366; wr31<=w_3_367; wr32<=w_3_368; wr33<=w_3_369; wr34<=w_3_370; wr35<=w_3_371; wr36<=w_3_372; wr37<=w_3_373; wr38<=w_3_374; wr39<=w_3_375; wr40<=w_3_376; wr41<=w_3_377; wr42<=w_3_378; wr43<=w_3_379; wr44<=w_3_380; wr45<=w_3_381; wr46<=w_3_382; wr47<=w_3_383; wr48<=w_3_384; wr49<=w_3_385; wr50<=w_3_386; wr51<=w_3_387; wr52<=w_3_388; wr53<=w_3_389; wr54<=w_3_390; wr55<=w_3_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd53:
					begin
						wr0<=w_3_392; wr1<=w_3_393; wr2<=w_3_394; wr3<=w_3_395; wr4<=w_3_396; wr5<=w_3_397; wr6<=w_3_398; wr7<=w_3_399; wr8<=w_3_400; wr9<=w_3_401; wr10<=w_3_402; wr11<=w_3_403; wr12<=w_3_404; wr13<=w_3_405; wr14<=w_3_406; wr15<=w_3_407; wr16<=w_3_408; wr17<=w_3_409; wr18<=w_3_410; wr19<=w_3_411; wr20<=w_3_412; wr21<=w_3_413; wr22<=w_3_414; wr23<=w_3_415; wr24<=w_3_416; wr25<=w_3_417; wr26<=w_3_418; wr27<=w_3_419; wr28<=w_3_420; wr29<=w_3_421; wr30<=w_3_422; wr31<=w_3_423; wr32<=w_3_424; wr33<=w_3_425; wr34<=w_3_426; wr35<=w_3_427; wr36<=w_3_428; wr37<=w_3_429; wr38<=w_3_430; wr39<=w_3_431; wr40<=w_3_432; wr41<=w_3_433; wr42<=w_3_434; wr43<=w_3_435; wr44<=w_3_436; wr45<=w_3_437; wr46<=w_3_438; wr47<=w_3_439; wr48<=w_3_440; wr49<=w_3_441; wr50<=w_3_442; wr51<=w_3_443; wr52<=w_3_444; wr53<=w_3_445; wr54<=w_3_446; wr55<=w_3_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd54:
					begin
						wr0<=w_3_448; wr1<=w_3_449; wr2<=w_3_450; wr3<=w_3_451; wr4<=w_3_452; wr5<=w_3_453; wr6<=w_3_454; wr7<=w_3_455; wr8<=w_3_456; wr9<=w_3_457; wr10<=w_3_458; wr11<=w_3_459; wr12<=w_3_460; wr13<=w_3_461; wr14<=w_3_462; wr15<=w_3_463; wr16<=w_3_464; wr17<=w_3_465; wr18<=w_3_466; wr19<=w_3_467; wr20<=w_3_468; wr21<=w_3_469; wr22<=w_3_470; wr23<=w_3_471; wr24<=w_3_472; wr25<=w_3_473; wr26<=w_3_474; wr27<=w_3_475; wr28<=w_3_476; wr29<=w_3_477; wr30<=w_3_478; wr31<=w_3_479; wr32<=w_3_480; wr33<=w_3_481; wr34<=w_3_482; wr35<=w_3_483; wr36<=w_3_484; wr37<=w_3_485; wr38<=w_3_486; wr39<=w_3_487; wr40<=w_3_488; wr41<=w_3_489; wr42<=w_3_490; wr43<=w_3_491; wr44<=w_3_492; wr45<=w_3_493; wr46<=w_3_494; wr47<=w_3_495; wr48<=w_3_496; wr49<=w_3_497; wr50<=w_3_498; wr51<=w_3_499; wr52<=w_3_500; wr53<=w_3_501; wr54<=w_3_502; wr55<=w_3_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd55:
					begin
						wr0<=w_3_504; wr1<=w_3_505; wr2<=w_3_506; wr3<=w_3_507; wr4<=w_3_508; wr5<=w_3_509; wr6<=w_3_510; wr7<=w_3_511; wr8<=w_3_512; wr9<=w_3_513; wr10<=w_3_514; wr11<=w_3_515; wr12<=w_3_516; wr13<=w_3_517; wr14<=w_3_518; wr15<=w_3_519; wr16<=w_3_520; wr17<=w_3_521; wr18<=w_3_522; wr19<=w_3_523; wr20<=w_3_524; wr21<=w_3_525; wr22<=w_3_526; wr23<=w_3_527; wr24<=w_3_528; wr25<=w_3_529; wr26<=w_3_530; wr27<=w_3_531; wr28<=w_3_532; wr29<=w_3_533; wr30<=w_3_534; wr31<=w_3_535; wr32<=w_3_536; wr33<=w_3_537; wr34<=w_3_538; wr35<=w_3_539; wr36<=w_3_540; wr37<=w_3_541; wr38<=w_3_542; wr39<=w_3_543; wr40<=w_3_544; wr41<=w_3_545; wr42<=w_3_546; wr43<=w_3_547; wr44<=w_3_548; wr45<=w_3_549; wr46<=w_3_550; wr47<=w_3_551; wr48<=w_3_552; wr49<=w_3_553; wr50<=w_3_554; wr51<=w_3_555; wr52<=w_3_556; wr53<=w_3_557; wr54<=w_3_558; wr55<=w_3_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd56:
					begin
						wr0<=w_3_560; wr1<=w_3_561; wr2<=w_3_562; wr3<=w_3_563; wr4<=w_3_564; wr5<=w_3_565; wr6<=w_3_566; wr7<=w_3_567; wr8<=w_3_568; wr9<=w_3_569; wr10<=w_3_570; wr11<=w_3_571; wr12<=w_3_572; wr13<=w_3_573; wr14<=w_3_574; wr15<=w_3_575; wr16<=w_3_576; wr17<=w_3_577; wr18<=w_3_578; wr19<=w_3_579; wr20<=w_3_580; wr21<=w_3_581; wr22<=w_3_582; wr23<=w_3_583; wr24<=w_3_584; wr25<=w_3_585; wr26<=w_3_586; wr27<=w_3_587; wr28<=w_3_588; wr29<=w_3_589; wr30<=w_3_590; wr31<=w_3_591; wr32<=w_3_592; wr33<=w_3_593; wr34<=w_3_594; wr35<=w_3_595; wr36<=w_3_596; wr37<=w_3_597; wr38<=w_3_598; wr39<=w_3_599; wr40<=w_3_600; wr41<=w_3_601; wr42<=w_3_602; wr43<=w_3_603; wr44<=w_3_604; wr45<=w_3_605; wr46<=w_3_606; wr47<=w_3_607; wr48<=w_3_608; wr49<=w_3_609; wr50<=w_3_610; wr51<=w_3_611; wr52<=w_3_612; wr53<=w_3_613; wr54<=w_3_614; wr55<=w_3_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd57:
					begin
						wr0<=w_3_616; wr1<=w_3_617; wr2<=w_3_618; wr3<=w_3_619; wr4<=w_3_620; wr5<=w_3_621; wr6<=w_3_622; wr7<=w_3_623; wr8<=w_3_624; wr9<=w_3_625; wr10<=w_3_626; wr11<=w_3_627; wr12<=w_3_628; wr13<=w_3_629; wr14<=w_3_630; wr15<=w_3_631; wr16<=w_3_632; wr17<=w_3_633; wr18<=w_3_634; wr19<=w_3_635; wr20<=w_3_636; wr21<=w_3_637; wr22<=w_3_638; wr23<=w_3_639; wr24<=w_3_640; wr25<=w_3_641; wr26<=w_3_642; wr27<=w_3_643; wr28<=w_3_644; wr29<=w_3_645; wr30<=w_3_646; wr31<=w_3_647; wr32<=w_3_648; wr33<=w_3_649; wr34<=w_3_650; wr35<=w_3_651; wr36<=w_3_652; wr37<=w_3_653; wr38<=w_3_654; wr39<=w_3_655; wr40<=w_3_656; wr41<=w_3_657; wr42<=w_3_658; wr43<=w_3_659; wr44<=w_3_660; wr45<=w_3_661; wr46<=w_3_662; wr47<=w_3_663; wr48<=w_3_664; wr49<=w_3_665; wr50<=w_3_666; wr51<=w_3_667; wr52<=w_3_668; wr53<=w_3_669; wr54<=w_3_670; wr55<=w_3_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd58:
					begin
						wr0<=w_3_672; wr1<=w_3_673; wr2<=w_3_674; wr3<=w_3_675; wr4<=w_3_676; wr5<=w_3_677; wr6<=w_3_678; wr7<=w_3_679; wr8<=w_3_680; wr9<=w_3_681; wr10<=w_3_682; wr11<=w_3_683; wr12<=w_3_684; wr13<=w_3_685; wr14<=w_3_686; wr15<=w_3_687; wr16<=w_3_688; wr17<=w_3_689; wr18<=w_3_690; wr19<=w_3_691; wr20<=w_3_692; wr21<=w_3_693; wr22<=w_3_694; wr23<=w_3_695; wr24<=w_3_696; wr25<=w_3_697; wr26<=w_3_698; wr27<=w_3_699; wr28<=w_3_700; wr29<=w_3_701; wr30<=w_3_702; wr31<=w_3_703; wr32<=w_3_704; wr33<=w_3_705; wr34<=w_3_706; wr35<=w_3_707; wr36<=w_3_708; wr37<=w_3_709; wr38<=w_3_710; wr39<=w_3_711; wr40<=w_3_712; wr41<=w_3_713; wr42<=w_3_714; wr43<=w_3_715; wr44<=w_3_716; wr45<=w_3_717; wr46<=w_3_718; wr47<=w_3_719; wr48<=w_3_720; wr49<=w_3_721; wr50<=w_3_722; wr51<=w_3_723; wr52<=w_3_724; wr53<=w_3_725; wr54<=w_3_726; wr55<=w_3_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd59:
					begin
						wr0<=w_3_728; wr1<=w_3_729; wr2<=w_3_730; wr3<=w_3_731; wr4<=w_3_732; wr5<=w_3_733; wr6<=w_3_734; wr7<=w_3_735; wr8<=w_3_736; wr9<=w_3_737; wr10<=w_3_738; wr11<=w_3_739; wr12<=w_3_740; wr13<=w_3_741; wr14<=w_3_742; wr15<=w_3_743; wr16<=w_3_744; wr17<=w_3_745; wr18<=w_3_746; wr19<=w_3_747; wr20<=w_3_748; wr21<=w_3_749; wr22<=w_3_750; wr23<=w_3_751; wr24<=w_3_752; wr25<=w_3_753; wr26<=w_3_754; wr27<=w_3_755; wr28<=w_3_756; wr29<=w_3_757; wr30<=w_3_758; wr31<=w_3_759; wr32<=w_3_760; wr33<=w_3_761; wr34<=w_3_762; wr35<=w_3_763; wr36<=w_3_764; wr37<=w_3_765; wr38<=w_3_766; wr39<=w_3_767; wr40<=w_3_768; wr41<=w_3_769; wr42<=w_3_770; wr43<=w_3_771; wr44<=w_3_772; wr45<=w_3_773; wr46<=w_3_774; wr47<=w_3_775; wr48<=w_3_776; wr49<=w_3_777; wr50<=w_3_778; wr51<=w_3_779; wr52<=w_3_780; wr53<=w_3_781; wr54<=w_3_782; wr55<=w_3_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd60:
					begin
						bias_p<=px_784;
						bias_w<=w_3_784;
						select<=select+1;
					end
				8'd61:
					begin
						wr0<=w_4_0; wr1<=w_4_1; wr2<=w_4_2; wr3<=w_4_3; wr4<=w_4_4; wr5<=w_4_5; wr6<=w_4_6; wr7<=w_4_7; wr8<=w_4_8; wr9<=w_4_9; wr10<=w_4_10; wr11<=w_4_11; wr12<=w_4_12; wr13<=w_4_13; wr14<=w_4_14; wr15<=w_4_15; wr16<=w_4_16; wr17<=w_4_17; wr18<=w_4_18; wr19<=w_4_19; wr20<=w_4_20; wr21<=w_4_21; wr22<=w_4_22; wr23<=w_4_23; wr24<=w_4_24; wr25<=w_4_25; wr26<=w_4_26; wr27<=w_4_27; wr28<=w_4_28; wr29<=w_4_29; wr30<=w_4_30; wr31<=w_4_31; wr32<=w_4_32; wr33<=w_4_33; wr34<=w_4_34; wr35<=w_4_35; wr36<=w_4_36; wr37<=w_4_37; wr38<=w_4_38; wr39<=w_4_39; wr40<=w_4_40; wr41<=w_4_41; wr42<=w_4_42; wr43<=w_4_43; wr44<=w_4_44; wr45<=w_4_45; wr46<=w_4_46; wr47<=w_4_47; wr48<=w_4_48; wr49<=w_4_49; wr50<=w_4_50; wr51<=w_4_51; wr52<=w_4_52; wr53<=w_4_53; wr54<=w_4_54; wr55<=w_4_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd62:
					begin
						wr0<=w_4_56; wr1<=w_4_57; wr2<=w_4_58; wr3<=w_4_59; wr4<=w_4_60; wr5<=w_4_61; wr6<=w_4_62; wr7<=w_4_63; wr8<=w_4_64; wr9<=w_4_65; wr10<=w_4_66; wr11<=w_4_67; wr12<=w_4_68; wr13<=w_4_69; wr14<=w_4_70; wr15<=w_4_71; wr16<=w_4_72; wr17<=w_4_73; wr18<=w_4_74; wr19<=w_4_75; wr20<=w_4_76; wr21<=w_4_77; wr22<=w_4_78; wr23<=w_4_79; wr24<=w_4_80; wr25<=w_4_81; wr26<=w_4_82; wr27<=w_4_83; wr28<=w_4_84; wr29<=w_4_85; wr30<=w_4_86; wr31<=w_4_87; wr32<=w_4_88; wr33<=w_4_89; wr34<=w_4_90; wr35<=w_4_91; wr36<=w_4_92; wr37<=w_4_93; wr38<=w_4_94; wr39<=w_4_95; wr40<=w_4_96; wr41<=w_4_97; wr42<=w_4_98; wr43<=w_4_99; wr44<=w_4_100; wr45<=w_4_101; wr46<=w_4_102; wr47<=w_4_103; wr48<=w_4_104; wr49<=w_4_105; wr50<=w_4_106; wr51<=w_4_107; wr52<=w_4_108; wr53<=w_4_109; wr54<=w_4_110; wr55<=w_4_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd63:
					begin
						wr0<=w_4_112; wr1<=w_4_113; wr2<=w_4_114; wr3<=w_4_115; wr4<=w_4_116; wr5<=w_4_117; wr6<=w_4_118; wr7<=w_4_119; wr8<=w_4_120; wr9<=w_4_121; wr10<=w_4_122; wr11<=w_4_123; wr12<=w_4_124; wr13<=w_4_125; wr14<=w_4_126; wr15<=w_4_127; wr16<=w_4_128; wr17<=w_4_129; wr18<=w_4_130; wr19<=w_4_131; wr20<=w_4_132; wr21<=w_4_133; wr22<=w_4_134; wr23<=w_4_135; wr24<=w_4_136; wr25<=w_4_137; wr26<=w_4_138; wr27<=w_4_139; wr28<=w_4_140; wr29<=w_4_141; wr30<=w_4_142; wr31<=w_4_143; wr32<=w_4_144; wr33<=w_4_145; wr34<=w_4_146; wr35<=w_4_147; wr36<=w_4_148; wr37<=w_4_149; wr38<=w_4_150; wr39<=w_4_151; wr40<=w_4_152; wr41<=w_4_153; wr42<=w_4_154; wr43<=w_4_155; wr44<=w_4_156; wr45<=w_4_157; wr46<=w_4_158; wr47<=w_4_159; wr48<=w_4_160; wr49<=w_4_161; wr50<=w_4_162; wr51<=w_4_163; wr52<=w_4_164; wr53<=w_4_165; wr54<=w_4_166; wr55<=w_4_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd64:
					begin
						wr0<=w_4_168; wr1<=w_4_169; wr2<=w_4_170; wr3<=w_4_171; wr4<=w_4_172; wr5<=w_4_173; wr6<=w_4_174; wr7<=w_4_175; wr8<=w_4_176; wr9<=w_4_177; wr10<=w_4_178; wr11<=w_4_179; wr12<=w_4_180; wr13<=w_4_181; wr14<=w_4_182; wr15<=w_4_183; wr16<=w_4_184; wr17<=w_4_185; wr18<=w_4_186; wr19<=w_4_187; wr20<=w_4_188; wr21<=w_4_189; wr22<=w_4_190; wr23<=w_4_191; wr24<=w_4_192; wr25<=w_4_193; wr26<=w_4_194; wr27<=w_4_195; wr28<=w_4_196; wr29<=w_4_197; wr30<=w_4_198; wr31<=w_4_199; wr32<=w_4_200; wr33<=w_4_201; wr34<=w_4_202; wr35<=w_4_203; wr36<=w_4_204; wr37<=w_4_205; wr38<=w_4_206; wr39<=w_4_207; wr40<=w_4_208; wr41<=w_4_209; wr42<=w_4_210; wr43<=w_4_211; wr44<=w_4_212; wr45<=w_4_213; wr46<=w_4_214; wr47<=w_4_215; wr48<=w_4_216; wr49<=w_4_217; wr50<=w_4_218; wr51<=w_4_219; wr52<=w_4_220; wr53<=w_4_221; wr54<=w_4_222; wr55<=w_4_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd65:
					begin
						wr0<=w_4_224; wr1<=w_4_225; wr2<=w_4_226; wr3<=w_4_227; wr4<=w_4_228; wr5<=w_4_229; wr6<=w_4_230; wr7<=w_4_231; wr8<=w_4_232; wr9<=w_4_233; wr10<=w_4_234; wr11<=w_4_235; wr12<=w_4_236; wr13<=w_4_237; wr14<=w_4_238; wr15<=w_4_239; wr16<=w_4_240; wr17<=w_4_241; wr18<=w_4_242; wr19<=w_4_243; wr20<=w_4_244; wr21<=w_4_245; wr22<=w_4_246; wr23<=w_4_247; wr24<=w_4_248; wr25<=w_4_249; wr26<=w_4_250; wr27<=w_4_251; wr28<=w_4_252; wr29<=w_4_253; wr30<=w_4_254; wr31<=w_4_255; wr32<=w_4_256; wr33<=w_4_257; wr34<=w_4_258; wr35<=w_4_259; wr36<=w_4_260; wr37<=w_4_261; wr38<=w_4_262; wr39<=w_4_263; wr40<=w_4_264; wr41<=w_4_265; wr42<=w_4_266; wr43<=w_4_267; wr44<=w_4_268; wr45<=w_4_269; wr46<=w_4_270; wr47<=w_4_271; wr48<=w_4_272; wr49<=w_4_273; wr50<=w_4_274; wr51<=w_4_275; wr52<=w_4_276; wr53<=w_4_277; wr54<=w_4_278; wr55<=w_4_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd66:
					begin
						wr0<=w_4_280; wr1<=w_4_281; wr2<=w_4_282; wr3<=w_4_283; wr4<=w_4_284; wr5<=w_4_285; wr6<=w_4_286; wr7<=w_4_287; wr8<=w_4_288; wr9<=w_4_289; wr10<=w_4_290; wr11<=w_4_291; wr12<=w_4_292; wr13<=w_4_293; wr14<=w_4_294; wr15<=w_4_295; wr16<=w_4_296; wr17<=w_4_297; wr18<=w_4_298; wr19<=w_4_299; wr20<=w_4_300; wr21<=w_4_301; wr22<=w_4_302; wr23<=w_4_303; wr24<=w_4_304; wr25<=w_4_305; wr26<=w_4_306; wr27<=w_4_307; wr28<=w_4_308; wr29<=w_4_309; wr30<=w_4_310; wr31<=w_4_311; wr32<=w_4_312; wr33<=w_4_313; wr34<=w_4_314; wr35<=w_4_315; wr36<=w_4_316; wr37<=w_4_317; wr38<=w_4_318; wr39<=w_4_319; wr40<=w_4_320; wr41<=w_4_321; wr42<=w_4_322; wr43<=w_4_323; wr44<=w_4_324; wr45<=w_4_325; wr46<=w_4_326; wr47<=w_4_327; wr48<=w_4_328; wr49<=w_4_329; wr50<=w_4_330; wr51<=w_4_331; wr52<=w_4_332; wr53<=w_4_333; wr54<=w_4_334; wr55<=w_4_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd67:
					begin
						wr0<=w_4_336; wr1<=w_4_337; wr2<=w_4_338; wr3<=w_4_339; wr4<=w_4_340; wr5<=w_4_341; wr6<=w_4_342; wr7<=w_4_343; wr8<=w_4_344; wr9<=w_4_345; wr10<=w_4_346; wr11<=w_4_347; wr12<=w_4_348; wr13<=w_4_349; wr14<=w_4_350; wr15<=w_4_351; wr16<=w_4_352; wr17<=w_4_353; wr18<=w_4_354; wr19<=w_4_355; wr20<=w_4_356; wr21<=w_4_357; wr22<=w_4_358; wr23<=w_4_359; wr24<=w_4_360; wr25<=w_4_361; wr26<=w_4_362; wr27<=w_4_363; wr28<=w_4_364; wr29<=w_4_365; wr30<=w_4_366; wr31<=w_4_367; wr32<=w_4_368; wr33<=w_4_369; wr34<=w_4_370; wr35<=w_4_371; wr36<=w_4_372; wr37<=w_4_373; wr38<=w_4_374; wr39<=w_4_375; wr40<=w_4_376; wr41<=w_4_377; wr42<=w_4_378; wr43<=w_4_379; wr44<=w_4_380; wr45<=w_4_381; wr46<=w_4_382; wr47<=w_4_383; wr48<=w_4_384; wr49<=w_4_385; wr50<=w_4_386; wr51<=w_4_387; wr52<=w_4_388; wr53<=w_4_389; wr54<=w_4_390; wr55<=w_4_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd68:
					begin
						wr0<=w_4_392; wr1<=w_4_393; wr2<=w_4_394; wr3<=w_4_395; wr4<=w_4_396; wr5<=w_4_397; wr6<=w_4_398; wr7<=w_4_399; wr8<=w_4_400; wr9<=w_4_401; wr10<=w_4_402; wr11<=w_4_403; wr12<=w_4_404; wr13<=w_4_405; wr14<=w_4_406; wr15<=w_4_407; wr16<=w_4_408; wr17<=w_4_409; wr18<=w_4_410; wr19<=w_4_411; wr20<=w_4_412; wr21<=w_4_413; wr22<=w_4_414; wr23<=w_4_415; wr24<=w_4_416; wr25<=w_4_417; wr26<=w_4_418; wr27<=w_4_419; wr28<=w_4_420; wr29<=w_4_421; wr30<=w_4_422; wr31<=w_4_423; wr32<=w_4_424; wr33<=w_4_425; wr34<=w_4_426; wr35<=w_4_427; wr36<=w_4_428; wr37<=w_4_429; wr38<=w_4_430; wr39<=w_4_431; wr40<=w_4_432; wr41<=w_4_433; wr42<=w_4_434; wr43<=w_4_435; wr44<=w_4_436; wr45<=w_4_437; wr46<=w_4_438; wr47<=w_4_439; wr48<=w_4_440; wr49<=w_4_441; wr50<=w_4_442; wr51<=w_4_443; wr52<=w_4_444; wr53<=w_4_445; wr54<=w_4_446; wr55<=w_4_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd69:
					begin
						wr0<=w_4_448; wr1<=w_4_449; wr2<=w_4_450; wr3<=w_4_451; wr4<=w_4_452; wr5<=w_4_453; wr6<=w_4_454; wr7<=w_4_455; wr8<=w_4_456; wr9<=w_4_457; wr10<=w_4_458; wr11<=w_4_459; wr12<=w_4_460; wr13<=w_4_461; wr14<=w_4_462; wr15<=w_4_463; wr16<=w_4_464; wr17<=w_4_465; wr18<=w_4_466; wr19<=w_4_467; wr20<=w_4_468; wr21<=w_4_469; wr22<=w_4_470; wr23<=w_4_471; wr24<=w_4_472; wr25<=w_4_473; wr26<=w_4_474; wr27<=w_4_475; wr28<=w_4_476; wr29<=w_4_477; wr30<=w_4_478; wr31<=w_4_479; wr32<=w_4_480; wr33<=w_4_481; wr34<=w_4_482; wr35<=w_4_483; wr36<=w_4_484; wr37<=w_4_485; wr38<=w_4_486; wr39<=w_4_487; wr40<=w_4_488; wr41<=w_4_489; wr42<=w_4_490; wr43<=w_4_491; wr44<=w_4_492; wr45<=w_4_493; wr46<=w_4_494; wr47<=w_4_495; wr48<=w_4_496; wr49<=w_4_497; wr50<=w_4_498; wr51<=w_4_499; wr52<=w_4_500; wr53<=w_4_501; wr54<=w_4_502; wr55<=w_4_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd70:
					begin
						wr0<=w_4_504; wr1<=w_4_505; wr2<=w_4_506; wr3<=w_4_507; wr4<=w_4_508; wr5<=w_4_509; wr6<=w_4_510; wr7<=w_4_511; wr8<=w_4_512; wr9<=w_4_513; wr10<=w_4_514; wr11<=w_4_515; wr12<=w_4_516; wr13<=w_4_517; wr14<=w_4_518; wr15<=w_4_519; wr16<=w_4_520; wr17<=w_4_521; wr18<=w_4_522; wr19<=w_4_523; wr20<=w_4_524; wr21<=w_4_525; wr22<=w_4_526; wr23<=w_4_527; wr24<=w_4_528; wr25<=w_4_529; wr26<=w_4_530; wr27<=w_4_531; wr28<=w_4_532; wr29<=w_4_533; wr30<=w_4_534; wr31<=w_4_535; wr32<=w_4_536; wr33<=w_4_537; wr34<=w_4_538; wr35<=w_4_539; wr36<=w_4_540; wr37<=w_4_541; wr38<=w_4_542; wr39<=w_4_543; wr40<=w_4_544; wr41<=w_4_545; wr42<=w_4_546; wr43<=w_4_547; wr44<=w_4_548; wr45<=w_4_549; wr46<=w_4_550; wr47<=w_4_551; wr48<=w_4_552; wr49<=w_4_553; wr50<=w_4_554; wr51<=w_4_555; wr52<=w_4_556; wr53<=w_4_557; wr54<=w_4_558; wr55<=w_4_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd71:
					begin
						wr0<=w_4_560; wr1<=w_4_561; wr2<=w_4_562; wr3<=w_4_563; wr4<=w_4_564; wr5<=w_4_565; wr6<=w_4_566; wr7<=w_4_567; wr8<=w_4_568; wr9<=w_4_569; wr10<=w_4_570; wr11<=w_4_571; wr12<=w_4_572; wr13<=w_4_573; wr14<=w_4_574; wr15<=w_4_575; wr16<=w_4_576; wr17<=w_4_577; wr18<=w_4_578; wr19<=w_4_579; wr20<=w_4_580; wr21<=w_4_581; wr22<=w_4_582; wr23<=w_4_583; wr24<=w_4_584; wr25<=w_4_585; wr26<=w_4_586; wr27<=w_4_587; wr28<=w_4_588; wr29<=w_4_589; wr30<=w_4_590; wr31<=w_4_591; wr32<=w_4_592; wr33<=w_4_593; wr34<=w_4_594; wr35<=w_4_595; wr36<=w_4_596; wr37<=w_4_597; wr38<=w_4_598; wr39<=w_4_599; wr40<=w_4_600; wr41<=w_4_601; wr42<=w_4_602; wr43<=w_4_603; wr44<=w_4_604; wr45<=w_4_605; wr46<=w_4_606; wr47<=w_4_607; wr48<=w_4_608; wr49<=w_4_609; wr50<=w_4_610; wr51<=w_4_611; wr52<=w_4_612; wr53<=w_4_613; wr54<=w_4_614; wr55<=w_4_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd72:
					begin
						wr0<=w_4_616; wr1<=w_4_617; wr2<=w_4_618; wr3<=w_4_619; wr4<=w_4_620; wr5<=w_4_621; wr6<=w_4_622; wr7<=w_4_623; wr8<=w_4_624; wr9<=w_4_625; wr10<=w_4_626; wr11<=w_4_627; wr12<=w_4_628; wr13<=w_4_629; wr14<=w_4_630; wr15<=w_4_631; wr16<=w_4_632; wr17<=w_4_633; wr18<=w_4_634; wr19<=w_4_635; wr20<=w_4_636; wr21<=w_4_637; wr22<=w_4_638; wr23<=w_4_639; wr24<=w_4_640; wr25<=w_4_641; wr26<=w_4_642; wr27<=w_4_643; wr28<=w_4_644; wr29<=w_4_645; wr30<=w_4_646; wr31<=w_4_647; wr32<=w_4_648; wr33<=w_4_649; wr34<=w_4_650; wr35<=w_4_651; wr36<=w_4_652; wr37<=w_4_653; wr38<=w_4_654; wr39<=w_4_655; wr40<=w_4_656; wr41<=w_4_657; wr42<=w_4_658; wr43<=w_4_659; wr44<=w_4_660; wr45<=w_4_661; wr46<=w_4_662; wr47<=w_4_663; wr48<=w_4_664; wr49<=w_4_665; wr50<=w_4_666; wr51<=w_4_667; wr52<=w_4_668; wr53<=w_4_669; wr54<=w_4_670; wr55<=w_4_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd73:
					begin
						wr0<=w_4_672; wr1<=w_4_673; wr2<=w_4_674; wr3<=w_4_675; wr4<=w_4_676; wr5<=w_4_677; wr6<=w_4_678; wr7<=w_4_679; wr8<=w_4_680; wr9<=w_4_681; wr10<=w_4_682; wr11<=w_4_683; wr12<=w_4_684; wr13<=w_4_685; wr14<=w_4_686; wr15<=w_4_687; wr16<=w_4_688; wr17<=w_4_689; wr18<=w_4_690; wr19<=w_4_691; wr20<=w_4_692; wr21<=w_4_693; wr22<=w_4_694; wr23<=w_4_695; wr24<=w_4_696; wr25<=w_4_697; wr26<=w_4_698; wr27<=w_4_699; wr28<=w_4_700; wr29<=w_4_701; wr30<=w_4_702; wr31<=w_4_703; wr32<=w_4_704; wr33<=w_4_705; wr34<=w_4_706; wr35<=w_4_707; wr36<=w_4_708; wr37<=w_4_709; wr38<=w_4_710; wr39<=w_4_711; wr40<=w_4_712; wr41<=w_4_713; wr42<=w_4_714; wr43<=w_4_715; wr44<=w_4_716; wr45<=w_4_717; wr46<=w_4_718; wr47<=w_4_719; wr48<=w_4_720; wr49<=w_4_721; wr50<=w_4_722; wr51<=w_4_723; wr52<=w_4_724; wr53<=w_4_725; wr54<=w_4_726; wr55<=w_4_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd74:
					begin
						wr0<=w_4_728; wr1<=w_4_729; wr2<=w_4_730; wr3<=w_4_731; wr4<=w_4_732; wr5<=w_4_733; wr6<=w_4_734; wr7<=w_4_735; wr8<=w_4_736; wr9<=w_4_737; wr10<=w_4_738; wr11<=w_4_739; wr12<=w_4_740; wr13<=w_4_741; wr14<=w_4_742; wr15<=w_4_743; wr16<=w_4_744; wr17<=w_4_745; wr18<=w_4_746; wr19<=w_4_747; wr20<=w_4_748; wr21<=w_4_749; wr22<=w_4_750; wr23<=w_4_751; wr24<=w_4_752; wr25<=w_4_753; wr26<=w_4_754; wr27<=w_4_755; wr28<=w_4_756; wr29<=w_4_757; wr30<=w_4_758; wr31<=w_4_759; wr32<=w_4_760; wr33<=w_4_761; wr34<=w_4_762; wr35<=w_4_763; wr36<=w_4_764; wr37<=w_4_765; wr38<=w_4_766; wr39<=w_4_767; wr40<=w_4_768; wr41<=w_4_769; wr42<=w_4_770; wr43<=w_4_771; wr44<=w_4_772; wr45<=w_4_773; wr46<=w_4_774; wr47<=w_4_775; wr48<=w_4_776; wr49<=w_4_777; wr50<=w_4_778; wr51<=w_4_779; wr52<=w_4_780; wr53<=w_4_781; wr54<=w_4_782; wr55<=w_4_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd75:
					begin
						bias_p<=px_784;
						bias_w<=w_4_784;
						select<=select+1;
					end
				8'd76:
					begin
						wr0<=w_5_0; wr1<=w_5_1; wr2<=w_5_2; wr3<=w_5_3; wr4<=w_5_4; wr5<=w_5_5; wr6<=w_5_6; wr7<=w_5_7; wr8<=w_5_8; wr9<=w_5_9; wr10<=w_5_10; wr11<=w_5_11; wr12<=w_5_12; wr13<=w_5_13; wr14<=w_5_14; wr15<=w_5_15; wr16<=w_5_16; wr17<=w_5_17; wr18<=w_5_18; wr19<=w_5_19; wr20<=w_5_20; wr21<=w_5_21; wr22<=w_5_22; wr23<=w_5_23; wr24<=w_5_24; wr25<=w_5_25; wr26<=w_5_26; wr27<=w_5_27; wr28<=w_5_28; wr29<=w_5_29; wr30<=w_5_30; wr31<=w_5_31; wr32<=w_5_32; wr33<=w_5_33; wr34<=w_5_34; wr35<=w_5_35; wr36<=w_5_36; wr37<=w_5_37; wr38<=w_5_38; wr39<=w_5_39; wr40<=w_5_40; wr41<=w_5_41; wr42<=w_5_42; wr43<=w_5_43; wr44<=w_5_44; wr45<=w_5_45; wr46<=w_5_46; wr47<=w_5_47; wr48<=w_5_48; wr49<=w_5_49; wr50<=w_5_50; wr51<=w_5_51; wr52<=w_5_52; wr53<=w_5_53; wr54<=w_5_54; wr55<=w_5_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd77:
					begin
						wr0<=w_5_56; wr1<=w_5_57; wr2<=w_5_58; wr3<=w_5_59; wr4<=w_5_60; wr5<=w_5_61; wr6<=w_5_62; wr7<=w_5_63; wr8<=w_5_64; wr9<=w_5_65; wr10<=w_5_66; wr11<=w_5_67; wr12<=w_5_68; wr13<=w_5_69; wr14<=w_5_70; wr15<=w_5_71; wr16<=w_5_72; wr17<=w_5_73; wr18<=w_5_74; wr19<=w_5_75; wr20<=w_5_76; wr21<=w_5_77; wr22<=w_5_78; wr23<=w_5_79; wr24<=w_5_80; wr25<=w_5_81; wr26<=w_5_82; wr27<=w_5_83; wr28<=w_5_84; wr29<=w_5_85; wr30<=w_5_86; wr31<=w_5_87; wr32<=w_5_88; wr33<=w_5_89; wr34<=w_5_90; wr35<=w_5_91; wr36<=w_5_92; wr37<=w_5_93; wr38<=w_5_94; wr39<=w_5_95; wr40<=w_5_96; wr41<=w_5_97; wr42<=w_5_98; wr43<=w_5_99; wr44<=w_5_100; wr45<=w_5_101; wr46<=w_5_102; wr47<=w_5_103; wr48<=w_5_104; wr49<=w_5_105; wr50<=w_5_106; wr51<=w_5_107; wr52<=w_5_108; wr53<=w_5_109; wr54<=w_5_110; wr55<=w_5_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd78:
					begin
						wr0<=w_5_112; wr1<=w_5_113; wr2<=w_5_114; wr3<=w_5_115; wr4<=w_5_116; wr5<=w_5_117; wr6<=w_5_118; wr7<=w_5_119; wr8<=w_5_120; wr9<=w_5_121; wr10<=w_5_122; wr11<=w_5_123; wr12<=w_5_124; wr13<=w_5_125; wr14<=w_5_126; wr15<=w_5_127; wr16<=w_5_128; wr17<=w_5_129; wr18<=w_5_130; wr19<=w_5_131; wr20<=w_5_132; wr21<=w_5_133; wr22<=w_5_134; wr23<=w_5_135; wr24<=w_5_136; wr25<=w_5_137; wr26<=w_5_138; wr27<=w_5_139; wr28<=w_5_140; wr29<=w_5_141; wr30<=w_5_142; wr31<=w_5_143; wr32<=w_5_144; wr33<=w_5_145; wr34<=w_5_146; wr35<=w_5_147; wr36<=w_5_148; wr37<=w_5_149; wr38<=w_5_150; wr39<=w_5_151; wr40<=w_5_152; wr41<=w_5_153; wr42<=w_5_154; wr43<=w_5_155; wr44<=w_5_156; wr45<=w_5_157; wr46<=w_5_158; wr47<=w_5_159; wr48<=w_5_160; wr49<=w_5_161; wr50<=w_5_162; wr51<=w_5_163; wr52<=w_5_164; wr53<=w_5_165; wr54<=w_5_166; wr55<=w_5_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd79:
					begin
						wr0<=w_5_168; wr1<=w_5_169; wr2<=w_5_170; wr3<=w_5_171; wr4<=w_5_172; wr5<=w_5_173; wr6<=w_5_174; wr7<=w_5_175; wr8<=w_5_176; wr9<=w_5_177; wr10<=w_5_178; wr11<=w_5_179; wr12<=w_5_180; wr13<=w_5_181; wr14<=w_5_182; wr15<=w_5_183; wr16<=w_5_184; wr17<=w_5_185; wr18<=w_5_186; wr19<=w_5_187; wr20<=w_5_188; wr21<=w_5_189; wr22<=w_5_190; wr23<=w_5_191; wr24<=w_5_192; wr25<=w_5_193; wr26<=w_5_194; wr27<=w_5_195; wr28<=w_5_196; wr29<=w_5_197; wr30<=w_5_198; wr31<=w_5_199; wr32<=w_5_200; wr33<=w_5_201; wr34<=w_5_202; wr35<=w_5_203; wr36<=w_5_204; wr37<=w_5_205; wr38<=w_5_206; wr39<=w_5_207; wr40<=w_5_208; wr41<=w_5_209; wr42<=w_5_210; wr43<=w_5_211; wr44<=w_5_212; wr45<=w_5_213; wr46<=w_5_214; wr47<=w_5_215; wr48<=w_5_216; wr49<=w_5_217; wr50<=w_5_218; wr51<=w_5_219; wr52<=w_5_220; wr53<=w_5_221; wr54<=w_5_222; wr55<=w_5_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd80:
					begin
						wr0<=w_5_224; wr1<=w_5_225; wr2<=w_5_226; wr3<=w_5_227; wr4<=w_5_228; wr5<=w_5_229; wr6<=w_5_230; wr7<=w_5_231; wr8<=w_5_232; wr9<=w_5_233; wr10<=w_5_234; wr11<=w_5_235; wr12<=w_5_236; wr13<=w_5_237; wr14<=w_5_238; wr15<=w_5_239; wr16<=w_5_240; wr17<=w_5_241; wr18<=w_5_242; wr19<=w_5_243; wr20<=w_5_244; wr21<=w_5_245; wr22<=w_5_246; wr23<=w_5_247; wr24<=w_5_248; wr25<=w_5_249; wr26<=w_5_250; wr27<=w_5_251; wr28<=w_5_252; wr29<=w_5_253; wr30<=w_5_254; wr31<=w_5_255; wr32<=w_5_256; wr33<=w_5_257; wr34<=w_5_258; wr35<=w_5_259; wr36<=w_5_260; wr37<=w_5_261; wr38<=w_5_262; wr39<=w_5_263; wr40<=w_5_264; wr41<=w_5_265; wr42<=w_5_266; wr43<=w_5_267; wr44<=w_5_268; wr45<=w_5_269; wr46<=w_5_270; wr47<=w_5_271; wr48<=w_5_272; wr49<=w_5_273; wr50<=w_5_274; wr51<=w_5_275; wr52<=w_5_276; wr53<=w_5_277; wr54<=w_5_278; wr55<=w_5_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd81:
					begin
						wr0<=w_5_280; wr1<=w_5_281; wr2<=w_5_282; wr3<=w_5_283; wr4<=w_5_284; wr5<=w_5_285; wr6<=w_5_286; wr7<=w_5_287; wr8<=w_5_288; wr9<=w_5_289; wr10<=w_5_290; wr11<=w_5_291; wr12<=w_5_292; wr13<=w_5_293; wr14<=w_5_294; wr15<=w_5_295; wr16<=w_5_296; wr17<=w_5_297; wr18<=w_5_298; wr19<=w_5_299; wr20<=w_5_300; wr21<=w_5_301; wr22<=w_5_302; wr23<=w_5_303; wr24<=w_5_304; wr25<=w_5_305; wr26<=w_5_306; wr27<=w_5_307; wr28<=w_5_308; wr29<=w_5_309; wr30<=w_5_310; wr31<=w_5_311; wr32<=w_5_312; wr33<=w_5_313; wr34<=w_5_314; wr35<=w_5_315; wr36<=w_5_316; wr37<=w_5_317; wr38<=w_5_318; wr39<=w_5_319; wr40<=w_5_320; wr41<=w_5_321; wr42<=w_5_322; wr43<=w_5_323; wr44<=w_5_324; wr45<=w_5_325; wr46<=w_5_326; wr47<=w_5_327; wr48<=w_5_328; wr49<=w_5_329; wr50<=w_5_330; wr51<=w_5_331; wr52<=w_5_332; wr53<=w_5_333; wr54<=w_5_334; wr55<=w_5_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd82:
					begin
						wr0<=w_5_336; wr1<=w_5_337; wr2<=w_5_338; wr3<=w_5_339; wr4<=w_5_340; wr5<=w_5_341; wr6<=w_5_342; wr7<=w_5_343; wr8<=w_5_344; wr9<=w_5_345; wr10<=w_5_346; wr11<=w_5_347; wr12<=w_5_348; wr13<=w_5_349; wr14<=w_5_350; wr15<=w_5_351; wr16<=w_5_352; wr17<=w_5_353; wr18<=w_5_354; wr19<=w_5_355; wr20<=w_5_356; wr21<=w_5_357; wr22<=w_5_358; wr23<=w_5_359; wr24<=w_5_360; wr25<=w_5_361; wr26<=w_5_362; wr27<=w_5_363; wr28<=w_5_364; wr29<=w_5_365; wr30<=w_5_366; wr31<=w_5_367; wr32<=w_5_368; wr33<=w_5_369; wr34<=w_5_370; wr35<=w_5_371; wr36<=w_5_372; wr37<=w_5_373; wr38<=w_5_374; wr39<=w_5_375; wr40<=w_5_376; wr41<=w_5_377; wr42<=w_5_378; wr43<=w_5_379; wr44<=w_5_380; wr45<=w_5_381; wr46<=w_5_382; wr47<=w_5_383; wr48<=w_5_384; wr49<=w_5_385; wr50<=w_5_386; wr51<=w_5_387; wr52<=w_5_388; wr53<=w_5_389; wr54<=w_5_390; wr55<=w_5_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd83:
					begin
						wr0<=w_5_392; wr1<=w_5_393; wr2<=w_5_394; wr3<=w_5_395; wr4<=w_5_396; wr5<=w_5_397; wr6<=w_5_398; wr7<=w_5_399; wr8<=w_5_400; wr9<=w_5_401; wr10<=w_5_402; wr11<=w_5_403; wr12<=w_5_404; wr13<=w_5_405; wr14<=w_5_406; wr15<=w_5_407; wr16<=w_5_408; wr17<=w_5_409; wr18<=w_5_410; wr19<=w_5_411; wr20<=w_5_412; wr21<=w_5_413; wr22<=w_5_414; wr23<=w_5_415; wr24<=w_5_416; wr25<=w_5_417; wr26<=w_5_418; wr27<=w_5_419; wr28<=w_5_420; wr29<=w_5_421; wr30<=w_5_422; wr31<=w_5_423; wr32<=w_5_424; wr33<=w_5_425; wr34<=w_5_426; wr35<=w_5_427; wr36<=w_5_428; wr37<=w_5_429; wr38<=w_5_430; wr39<=w_5_431; wr40<=w_5_432; wr41<=w_5_433; wr42<=w_5_434; wr43<=w_5_435; wr44<=w_5_436; wr45<=w_5_437; wr46<=w_5_438; wr47<=w_5_439; wr48<=w_5_440; wr49<=w_5_441; wr50<=w_5_442; wr51<=w_5_443; wr52<=w_5_444; wr53<=w_5_445; wr54<=w_5_446; wr55<=w_5_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd84:
					begin
						wr0<=w_5_448; wr1<=w_5_449; wr2<=w_5_450; wr3<=w_5_451; wr4<=w_5_452; wr5<=w_5_453; wr6<=w_5_454; wr7<=w_5_455; wr8<=w_5_456; wr9<=w_5_457; wr10<=w_5_458; wr11<=w_5_459; wr12<=w_5_460; wr13<=w_5_461; wr14<=w_5_462; wr15<=w_5_463; wr16<=w_5_464; wr17<=w_5_465; wr18<=w_5_466; wr19<=w_5_467; wr20<=w_5_468; wr21<=w_5_469; wr22<=w_5_470; wr23<=w_5_471; wr24<=w_5_472; wr25<=w_5_473; wr26<=w_5_474; wr27<=w_5_475; wr28<=w_5_476; wr29<=w_5_477; wr30<=w_5_478; wr31<=w_5_479; wr32<=w_5_480; wr33<=w_5_481; wr34<=w_5_482; wr35<=w_5_483; wr36<=w_5_484; wr37<=w_5_485; wr38<=w_5_486; wr39<=w_5_487; wr40<=w_5_488; wr41<=w_5_489; wr42<=w_5_490; wr43<=w_5_491; wr44<=w_5_492; wr45<=w_5_493; wr46<=w_5_494; wr47<=w_5_495; wr48<=w_5_496; wr49<=w_5_497; wr50<=w_5_498; wr51<=w_5_499; wr52<=w_5_500; wr53<=w_5_501; wr54<=w_5_502; wr55<=w_5_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd85:
					begin
						wr0<=w_5_504; wr1<=w_5_505; wr2<=w_5_506; wr3<=w_5_507; wr4<=w_5_508; wr5<=w_5_509; wr6<=w_5_510; wr7<=w_5_511; wr8<=w_5_512; wr9<=w_5_513; wr10<=w_5_514; wr11<=w_5_515; wr12<=w_5_516; wr13<=w_5_517; wr14<=w_5_518; wr15<=w_5_519; wr16<=w_5_520; wr17<=w_5_521; wr18<=w_5_522; wr19<=w_5_523; wr20<=w_5_524; wr21<=w_5_525; wr22<=w_5_526; wr23<=w_5_527; wr24<=w_5_528; wr25<=w_5_529; wr26<=w_5_530; wr27<=w_5_531; wr28<=w_5_532; wr29<=w_5_533; wr30<=w_5_534; wr31<=w_5_535; wr32<=w_5_536; wr33<=w_5_537; wr34<=w_5_538; wr35<=w_5_539; wr36<=w_5_540; wr37<=w_5_541; wr38<=w_5_542; wr39<=w_5_543; wr40<=w_5_544; wr41<=w_5_545; wr42<=w_5_546; wr43<=w_5_547; wr44<=w_5_548; wr45<=w_5_549; wr46<=w_5_550; wr47<=w_5_551; wr48<=w_5_552; wr49<=w_5_553; wr50<=w_5_554; wr51<=w_5_555; wr52<=w_5_556; wr53<=w_5_557; wr54<=w_5_558; wr55<=w_5_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd86:
					begin
						wr0<=w_5_560; wr1<=w_5_561; wr2<=w_5_562; wr3<=w_5_563; wr4<=w_5_564; wr5<=w_5_565; wr6<=w_5_566; wr7<=w_5_567; wr8<=w_5_568; wr9<=w_5_569; wr10<=w_5_570; wr11<=w_5_571; wr12<=w_5_572; wr13<=w_5_573; wr14<=w_5_574; wr15<=w_5_575; wr16<=w_5_576; wr17<=w_5_577; wr18<=w_5_578; wr19<=w_5_579; wr20<=w_5_580; wr21<=w_5_581; wr22<=w_5_582; wr23<=w_5_583; wr24<=w_5_584; wr25<=w_5_585; wr26<=w_5_586; wr27<=w_5_587; wr28<=w_5_588; wr29<=w_5_589; wr30<=w_5_590; wr31<=w_5_591; wr32<=w_5_592; wr33<=w_5_593; wr34<=w_5_594; wr35<=w_5_595; wr36<=w_5_596; wr37<=w_5_597; wr38<=w_5_598; wr39<=w_5_599; wr40<=w_5_600; wr41<=w_5_601; wr42<=w_5_602; wr43<=w_5_603; wr44<=w_5_604; wr45<=w_5_605; wr46<=w_5_606; wr47<=w_5_607; wr48<=w_5_608; wr49<=w_5_609; wr50<=w_5_610; wr51<=w_5_611; wr52<=w_5_612; wr53<=w_5_613; wr54<=w_5_614; wr55<=w_5_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd87:
					begin
						wr0<=w_5_616; wr1<=w_5_617; wr2<=w_5_618; wr3<=w_5_619; wr4<=w_5_620; wr5<=w_5_621; wr6<=w_5_622; wr7<=w_5_623; wr8<=w_5_624; wr9<=w_5_625; wr10<=w_5_626; wr11<=w_5_627; wr12<=w_5_628; wr13<=w_5_629; wr14<=w_5_630; wr15<=w_5_631; wr16<=w_5_632; wr17<=w_5_633; wr18<=w_5_634; wr19<=w_5_635; wr20<=w_5_636; wr21<=w_5_637; wr22<=w_5_638; wr23<=w_5_639; wr24<=w_5_640; wr25<=w_5_641; wr26<=w_5_642; wr27<=w_5_643; wr28<=w_5_644; wr29<=w_5_645; wr30<=w_5_646; wr31<=w_5_647; wr32<=w_5_648; wr33<=w_5_649; wr34<=w_5_650; wr35<=w_5_651; wr36<=w_5_652; wr37<=w_5_653; wr38<=w_5_654; wr39<=w_5_655; wr40<=w_5_656; wr41<=w_5_657; wr42<=w_5_658; wr43<=w_5_659; wr44<=w_5_660; wr45<=w_5_661; wr46<=w_5_662; wr47<=w_5_663; wr48<=w_5_664; wr49<=w_5_665; wr50<=w_5_666; wr51<=w_5_667; wr52<=w_5_668; wr53<=w_5_669; wr54<=w_5_670; wr55<=w_5_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd88:
					begin
						wr0<=w_5_672; wr1<=w_5_673; wr2<=w_5_674; wr3<=w_5_675; wr4<=w_5_676; wr5<=w_5_677; wr6<=w_5_678; wr7<=w_5_679; wr8<=w_5_680; wr9<=w_5_681; wr10<=w_5_682; wr11<=w_5_683; wr12<=w_5_684; wr13<=w_5_685; wr14<=w_5_686; wr15<=w_5_687; wr16<=w_5_688; wr17<=w_5_689; wr18<=w_5_690; wr19<=w_5_691; wr20<=w_5_692; wr21<=w_5_693; wr22<=w_5_694; wr23<=w_5_695; wr24<=w_5_696; wr25<=w_5_697; wr26<=w_5_698; wr27<=w_5_699; wr28<=w_5_700; wr29<=w_5_701; wr30<=w_5_702; wr31<=w_5_703; wr32<=w_5_704; wr33<=w_5_705; wr34<=w_5_706; wr35<=w_5_707; wr36<=w_5_708; wr37<=w_5_709; wr38<=w_5_710; wr39<=w_5_711; wr40<=w_5_712; wr41<=w_5_713; wr42<=w_5_714; wr43<=w_5_715; wr44<=w_5_716; wr45<=w_5_717; wr46<=w_5_718; wr47<=w_5_719; wr48<=w_5_720; wr49<=w_5_721; wr50<=w_5_722; wr51<=w_5_723; wr52<=w_5_724; wr53<=w_5_725; wr54<=w_5_726; wr55<=w_5_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd89:
					begin
						wr0<=w_5_728; wr1<=w_5_729; wr2<=w_5_730; wr3<=w_5_731; wr4<=w_5_732; wr5<=w_5_733; wr6<=w_5_734; wr7<=w_5_735; wr8<=w_5_736; wr9<=w_5_737; wr10<=w_5_738; wr11<=w_5_739; wr12<=w_5_740; wr13<=w_5_741; wr14<=w_5_742; wr15<=w_5_743; wr16<=w_5_744; wr17<=w_5_745; wr18<=w_5_746; wr19<=w_5_747; wr20<=w_5_748; wr21<=w_5_749; wr22<=w_5_750; wr23<=w_5_751; wr24<=w_5_752; wr25<=w_5_753; wr26<=w_5_754; wr27<=w_5_755; wr28<=w_5_756; wr29<=w_5_757; wr30<=w_5_758; wr31<=w_5_759; wr32<=w_5_760; wr33<=w_5_761; wr34<=w_5_762; wr35<=w_5_763; wr36<=w_5_764; wr37<=w_5_765; wr38<=w_5_766; wr39<=w_5_767; wr40<=w_5_768; wr41<=w_5_769; wr42<=w_5_770; wr43<=w_5_771; wr44<=w_5_772; wr45<=w_5_773; wr46<=w_5_774; wr47<=w_5_775; wr48<=w_5_776; wr49<=w_5_777; wr50<=w_5_778; wr51<=w_5_779; wr52<=w_5_780; wr53<=w_5_781; wr54<=w_5_782; wr55<=w_5_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd90:
					begin
						bias_p<=px_784;
						bias_w<=w_5_784;
						select<=select+1;
					end
				8'd91:
					begin
						wr0<=w_6_0; wr1<=w_6_1; wr2<=w_6_2; wr3<=w_6_3; wr4<=w_6_4; wr5<=w_6_5; wr6<=w_6_6; wr7<=w_6_7; wr8<=w_6_8; wr9<=w_6_9; wr10<=w_6_10; wr11<=w_6_11; wr12<=w_6_12; wr13<=w_6_13; wr14<=w_6_14; wr15<=w_6_15; wr16<=w_6_16; wr17<=w_6_17; wr18<=w_6_18; wr19<=w_6_19; wr20<=w_6_20; wr21<=w_6_21; wr22<=w_6_22; wr23<=w_6_23; wr24<=w_6_24; wr25<=w_6_25; wr26<=w_6_26; wr27<=w_6_27; wr28<=w_6_28; wr29<=w_6_29; wr30<=w_6_30; wr31<=w_6_31; wr32<=w_6_32; wr33<=w_6_33; wr34<=w_6_34; wr35<=w_6_35; wr36<=w_6_36; wr37<=w_6_37; wr38<=w_6_38; wr39<=w_6_39; wr40<=w_6_40; wr41<=w_6_41; wr42<=w_6_42; wr43<=w_6_43; wr44<=w_6_44; wr45<=w_6_45; wr46<=w_6_46; wr47<=w_6_47; wr48<=w_6_48; wr49<=w_6_49; wr50<=w_6_50; wr51<=w_6_51; wr52<=w_6_52; wr53<=w_6_53; wr54<=w_6_54; wr55<=w_6_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd92:
					begin
						wr0<=w_6_56; wr1<=w_6_57; wr2<=w_6_58; wr3<=w_6_59; wr4<=w_6_60; wr5<=w_6_61; wr6<=w_6_62; wr7<=w_6_63; wr8<=w_6_64; wr9<=w_6_65; wr10<=w_6_66; wr11<=w_6_67; wr12<=w_6_68; wr13<=w_6_69; wr14<=w_6_70; wr15<=w_6_71; wr16<=w_6_72; wr17<=w_6_73; wr18<=w_6_74; wr19<=w_6_75; wr20<=w_6_76; wr21<=w_6_77; wr22<=w_6_78; wr23<=w_6_79; wr24<=w_6_80; wr25<=w_6_81; wr26<=w_6_82; wr27<=w_6_83; wr28<=w_6_84; wr29<=w_6_85; wr30<=w_6_86; wr31<=w_6_87; wr32<=w_6_88; wr33<=w_6_89; wr34<=w_6_90; wr35<=w_6_91; wr36<=w_6_92; wr37<=w_6_93; wr38<=w_6_94; wr39<=w_6_95; wr40<=w_6_96; wr41<=w_6_97; wr42<=w_6_98; wr43<=w_6_99; wr44<=w_6_100; wr45<=w_6_101; wr46<=w_6_102; wr47<=w_6_103; wr48<=w_6_104; wr49<=w_6_105; wr50<=w_6_106; wr51<=w_6_107; wr52<=w_6_108; wr53<=w_6_109; wr54<=w_6_110; wr55<=w_6_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd93:
					begin
						wr0<=w_6_112; wr1<=w_6_113; wr2<=w_6_114; wr3<=w_6_115; wr4<=w_6_116; wr5<=w_6_117; wr6<=w_6_118; wr7<=w_6_119; wr8<=w_6_120; wr9<=w_6_121; wr10<=w_6_122; wr11<=w_6_123; wr12<=w_6_124; wr13<=w_6_125; wr14<=w_6_126; wr15<=w_6_127; wr16<=w_6_128; wr17<=w_6_129; wr18<=w_6_130; wr19<=w_6_131; wr20<=w_6_132; wr21<=w_6_133; wr22<=w_6_134; wr23<=w_6_135; wr24<=w_6_136; wr25<=w_6_137; wr26<=w_6_138; wr27<=w_6_139; wr28<=w_6_140; wr29<=w_6_141; wr30<=w_6_142; wr31<=w_6_143; wr32<=w_6_144; wr33<=w_6_145; wr34<=w_6_146; wr35<=w_6_147; wr36<=w_6_148; wr37<=w_6_149; wr38<=w_6_150; wr39<=w_6_151; wr40<=w_6_152; wr41<=w_6_153; wr42<=w_6_154; wr43<=w_6_155; wr44<=w_6_156; wr45<=w_6_157; wr46<=w_6_158; wr47<=w_6_159; wr48<=w_6_160; wr49<=w_6_161; wr50<=w_6_162; wr51<=w_6_163; wr52<=w_6_164; wr53<=w_6_165; wr54<=w_6_166; wr55<=w_6_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd94:
					begin
						wr0<=w_6_168; wr1<=w_6_169; wr2<=w_6_170; wr3<=w_6_171; wr4<=w_6_172; wr5<=w_6_173; wr6<=w_6_174; wr7<=w_6_175; wr8<=w_6_176; wr9<=w_6_177; wr10<=w_6_178; wr11<=w_6_179; wr12<=w_6_180; wr13<=w_6_181; wr14<=w_6_182; wr15<=w_6_183; wr16<=w_6_184; wr17<=w_6_185; wr18<=w_6_186; wr19<=w_6_187; wr20<=w_6_188; wr21<=w_6_189; wr22<=w_6_190; wr23<=w_6_191; wr24<=w_6_192; wr25<=w_6_193; wr26<=w_6_194; wr27<=w_6_195; wr28<=w_6_196; wr29<=w_6_197; wr30<=w_6_198; wr31<=w_6_199; wr32<=w_6_200; wr33<=w_6_201; wr34<=w_6_202; wr35<=w_6_203; wr36<=w_6_204; wr37<=w_6_205; wr38<=w_6_206; wr39<=w_6_207; wr40<=w_6_208; wr41<=w_6_209; wr42<=w_6_210; wr43<=w_6_211; wr44<=w_6_212; wr45<=w_6_213; wr46<=w_6_214; wr47<=w_6_215; wr48<=w_6_216; wr49<=w_6_217; wr50<=w_6_218; wr51<=w_6_219; wr52<=w_6_220; wr53<=w_6_221; wr54<=w_6_222; wr55<=w_6_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd95:
					begin
						wr0<=w_6_224; wr1<=w_6_225; wr2<=w_6_226; wr3<=w_6_227; wr4<=w_6_228; wr5<=w_6_229; wr6<=w_6_230; wr7<=w_6_231; wr8<=w_6_232; wr9<=w_6_233; wr10<=w_6_234; wr11<=w_6_235; wr12<=w_6_236; wr13<=w_6_237; wr14<=w_6_238; wr15<=w_6_239; wr16<=w_6_240; wr17<=w_6_241; wr18<=w_6_242; wr19<=w_6_243; wr20<=w_6_244; wr21<=w_6_245; wr22<=w_6_246; wr23<=w_6_247; wr24<=w_6_248; wr25<=w_6_249; wr26<=w_6_250; wr27<=w_6_251; wr28<=w_6_252; wr29<=w_6_253; wr30<=w_6_254; wr31<=w_6_255; wr32<=w_6_256; wr33<=w_6_257; wr34<=w_6_258; wr35<=w_6_259; wr36<=w_6_260; wr37<=w_6_261; wr38<=w_6_262; wr39<=w_6_263; wr40<=w_6_264; wr41<=w_6_265; wr42<=w_6_266; wr43<=w_6_267; wr44<=w_6_268; wr45<=w_6_269; wr46<=w_6_270; wr47<=w_6_271; wr48<=w_6_272; wr49<=w_6_273; wr50<=w_6_274; wr51<=w_6_275; wr52<=w_6_276; wr53<=w_6_277; wr54<=w_6_278; wr55<=w_6_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd96:
					begin
						wr0<=w_6_280; wr1<=w_6_281; wr2<=w_6_282; wr3<=w_6_283; wr4<=w_6_284; wr5<=w_6_285; wr6<=w_6_286; wr7<=w_6_287; wr8<=w_6_288; wr9<=w_6_289; wr10<=w_6_290; wr11<=w_6_291; wr12<=w_6_292; wr13<=w_6_293; wr14<=w_6_294; wr15<=w_6_295; wr16<=w_6_296; wr17<=w_6_297; wr18<=w_6_298; wr19<=w_6_299; wr20<=w_6_300; wr21<=w_6_301; wr22<=w_6_302; wr23<=w_6_303; wr24<=w_6_304; wr25<=w_6_305; wr26<=w_6_306; wr27<=w_6_307; wr28<=w_6_308; wr29<=w_6_309; wr30<=w_6_310; wr31<=w_6_311; wr32<=w_6_312; wr33<=w_6_313; wr34<=w_6_314; wr35<=w_6_315; wr36<=w_6_316; wr37<=w_6_317; wr38<=w_6_318; wr39<=w_6_319; wr40<=w_6_320; wr41<=w_6_321; wr42<=w_6_322; wr43<=w_6_323; wr44<=w_6_324; wr45<=w_6_325; wr46<=w_6_326; wr47<=w_6_327; wr48<=w_6_328; wr49<=w_6_329; wr50<=w_6_330; wr51<=w_6_331; wr52<=w_6_332; wr53<=w_6_333; wr54<=w_6_334; wr55<=w_6_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd97:
					begin
						wr0<=w_6_336; wr1<=w_6_337; wr2<=w_6_338; wr3<=w_6_339; wr4<=w_6_340; wr5<=w_6_341; wr6<=w_6_342; wr7<=w_6_343; wr8<=w_6_344; wr9<=w_6_345; wr10<=w_6_346; wr11<=w_6_347; wr12<=w_6_348; wr13<=w_6_349; wr14<=w_6_350; wr15<=w_6_351; wr16<=w_6_352; wr17<=w_6_353; wr18<=w_6_354; wr19<=w_6_355; wr20<=w_6_356; wr21<=w_6_357; wr22<=w_6_358; wr23<=w_6_359; wr24<=w_6_360; wr25<=w_6_361; wr26<=w_6_362; wr27<=w_6_363; wr28<=w_6_364; wr29<=w_6_365; wr30<=w_6_366; wr31<=w_6_367; wr32<=w_6_368; wr33<=w_6_369; wr34<=w_6_370; wr35<=w_6_371; wr36<=w_6_372; wr37<=w_6_373; wr38<=w_6_374; wr39<=w_6_375; wr40<=w_6_376; wr41<=w_6_377; wr42<=w_6_378; wr43<=w_6_379; wr44<=w_6_380; wr45<=w_6_381; wr46<=w_6_382; wr47<=w_6_383; wr48<=w_6_384; wr49<=w_6_385; wr50<=w_6_386; wr51<=w_6_387; wr52<=w_6_388; wr53<=w_6_389; wr54<=w_6_390; wr55<=w_6_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd98:
					begin
						wr0<=w_6_392; wr1<=w_6_393; wr2<=w_6_394; wr3<=w_6_395; wr4<=w_6_396; wr5<=w_6_397; wr6<=w_6_398; wr7<=w_6_399; wr8<=w_6_400; wr9<=w_6_401; wr10<=w_6_402; wr11<=w_6_403; wr12<=w_6_404; wr13<=w_6_405; wr14<=w_6_406; wr15<=w_6_407; wr16<=w_6_408; wr17<=w_6_409; wr18<=w_6_410; wr19<=w_6_411; wr20<=w_6_412; wr21<=w_6_413; wr22<=w_6_414; wr23<=w_6_415; wr24<=w_6_416; wr25<=w_6_417; wr26<=w_6_418; wr27<=w_6_419; wr28<=w_6_420; wr29<=w_6_421; wr30<=w_6_422; wr31<=w_6_423; wr32<=w_6_424; wr33<=w_6_425; wr34<=w_6_426; wr35<=w_6_427; wr36<=w_6_428; wr37<=w_6_429; wr38<=w_6_430; wr39<=w_6_431; wr40<=w_6_432; wr41<=w_6_433; wr42<=w_6_434; wr43<=w_6_435; wr44<=w_6_436; wr45<=w_6_437; wr46<=w_6_438; wr47<=w_6_439; wr48<=w_6_440; wr49<=w_6_441; wr50<=w_6_442; wr51<=w_6_443; wr52<=w_6_444; wr53<=w_6_445; wr54<=w_6_446; wr55<=w_6_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd99:
					begin
						wr0<=w_6_448; wr1<=w_6_449; wr2<=w_6_450; wr3<=w_6_451; wr4<=w_6_452; wr5<=w_6_453; wr6<=w_6_454; wr7<=w_6_455; wr8<=w_6_456; wr9<=w_6_457; wr10<=w_6_458; wr11<=w_6_459; wr12<=w_6_460; wr13<=w_6_461; wr14<=w_6_462; wr15<=w_6_463; wr16<=w_6_464; wr17<=w_6_465; wr18<=w_6_466; wr19<=w_6_467; wr20<=w_6_468; wr21<=w_6_469; wr22<=w_6_470; wr23<=w_6_471; wr24<=w_6_472; wr25<=w_6_473; wr26<=w_6_474; wr27<=w_6_475; wr28<=w_6_476; wr29<=w_6_477; wr30<=w_6_478; wr31<=w_6_479; wr32<=w_6_480; wr33<=w_6_481; wr34<=w_6_482; wr35<=w_6_483; wr36<=w_6_484; wr37<=w_6_485; wr38<=w_6_486; wr39<=w_6_487; wr40<=w_6_488; wr41<=w_6_489; wr42<=w_6_490; wr43<=w_6_491; wr44<=w_6_492; wr45<=w_6_493; wr46<=w_6_494; wr47<=w_6_495; wr48<=w_6_496; wr49<=w_6_497; wr50<=w_6_498; wr51<=w_6_499; wr52<=w_6_500; wr53<=w_6_501; wr54<=w_6_502; wr55<=w_6_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd100:
					begin
						wr0<=w_6_504; wr1<=w_6_505; wr2<=w_6_506; wr3<=w_6_507; wr4<=w_6_508; wr5<=w_6_509; wr6<=w_6_510; wr7<=w_6_511; wr8<=w_6_512; wr9<=w_6_513; wr10<=w_6_514; wr11<=w_6_515; wr12<=w_6_516; wr13<=w_6_517; wr14<=w_6_518; wr15<=w_6_519; wr16<=w_6_520; wr17<=w_6_521; wr18<=w_6_522; wr19<=w_6_523; wr20<=w_6_524; wr21<=w_6_525; wr22<=w_6_526; wr23<=w_6_527; wr24<=w_6_528; wr25<=w_6_529; wr26<=w_6_530; wr27<=w_6_531; wr28<=w_6_532; wr29<=w_6_533; wr30<=w_6_534; wr31<=w_6_535; wr32<=w_6_536; wr33<=w_6_537; wr34<=w_6_538; wr35<=w_6_539; wr36<=w_6_540; wr37<=w_6_541; wr38<=w_6_542; wr39<=w_6_543; wr40<=w_6_544; wr41<=w_6_545; wr42<=w_6_546; wr43<=w_6_547; wr44<=w_6_548; wr45<=w_6_549; wr46<=w_6_550; wr47<=w_6_551; wr48<=w_6_552; wr49<=w_6_553; wr50<=w_6_554; wr51<=w_6_555; wr52<=w_6_556; wr53<=w_6_557; wr54<=w_6_558; wr55<=w_6_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd101:
					begin
						wr0<=w_6_560; wr1<=w_6_561; wr2<=w_6_562; wr3<=w_6_563; wr4<=w_6_564; wr5<=w_6_565; wr6<=w_6_566; wr7<=w_6_567; wr8<=w_6_568; wr9<=w_6_569; wr10<=w_6_570; wr11<=w_6_571; wr12<=w_6_572; wr13<=w_6_573; wr14<=w_6_574; wr15<=w_6_575; wr16<=w_6_576; wr17<=w_6_577; wr18<=w_6_578; wr19<=w_6_579; wr20<=w_6_580; wr21<=w_6_581; wr22<=w_6_582; wr23<=w_6_583; wr24<=w_6_584; wr25<=w_6_585; wr26<=w_6_586; wr27<=w_6_587; wr28<=w_6_588; wr29<=w_6_589; wr30<=w_6_590; wr31<=w_6_591; wr32<=w_6_592; wr33<=w_6_593; wr34<=w_6_594; wr35<=w_6_595; wr36<=w_6_596; wr37<=w_6_597; wr38<=w_6_598; wr39<=w_6_599; wr40<=w_6_600; wr41<=w_6_601; wr42<=w_6_602; wr43<=w_6_603; wr44<=w_6_604; wr45<=w_6_605; wr46<=w_6_606; wr47<=w_6_607; wr48<=w_6_608; wr49<=w_6_609; wr50<=w_6_610; wr51<=w_6_611; wr52<=w_6_612; wr53<=w_6_613; wr54<=w_6_614; wr55<=w_6_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd102:
					begin
						wr0<=w_6_616; wr1<=w_6_617; wr2<=w_6_618; wr3<=w_6_619; wr4<=w_6_620; wr5<=w_6_621; wr6<=w_6_622; wr7<=w_6_623; wr8<=w_6_624; wr9<=w_6_625; wr10<=w_6_626; wr11<=w_6_627; wr12<=w_6_628; wr13<=w_6_629; wr14<=w_6_630; wr15<=w_6_631; wr16<=w_6_632; wr17<=w_6_633; wr18<=w_6_634; wr19<=w_6_635; wr20<=w_6_636; wr21<=w_6_637; wr22<=w_6_638; wr23<=w_6_639; wr24<=w_6_640; wr25<=w_6_641; wr26<=w_6_642; wr27<=w_6_643; wr28<=w_6_644; wr29<=w_6_645; wr30<=w_6_646; wr31<=w_6_647; wr32<=w_6_648; wr33<=w_6_649; wr34<=w_6_650; wr35<=w_6_651; wr36<=w_6_652; wr37<=w_6_653; wr38<=w_6_654; wr39<=w_6_655; wr40<=w_6_656; wr41<=w_6_657; wr42<=w_6_658; wr43<=w_6_659; wr44<=w_6_660; wr45<=w_6_661; wr46<=w_6_662; wr47<=w_6_663; wr48<=w_6_664; wr49<=w_6_665; wr50<=w_6_666; wr51<=w_6_667; wr52<=w_6_668; wr53<=w_6_669; wr54<=w_6_670; wr55<=w_6_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd103:
					begin
						wr0<=w_6_672; wr1<=w_6_673; wr2<=w_6_674; wr3<=w_6_675; wr4<=w_6_676; wr5<=w_6_677; wr6<=w_6_678; wr7<=w_6_679; wr8<=w_6_680; wr9<=w_6_681; wr10<=w_6_682; wr11<=w_6_683; wr12<=w_6_684; wr13<=w_6_685; wr14<=w_6_686; wr15<=w_6_687; wr16<=w_6_688; wr17<=w_6_689; wr18<=w_6_690; wr19<=w_6_691; wr20<=w_6_692; wr21<=w_6_693; wr22<=w_6_694; wr23<=w_6_695; wr24<=w_6_696; wr25<=w_6_697; wr26<=w_6_698; wr27<=w_6_699; wr28<=w_6_700; wr29<=w_6_701; wr30<=w_6_702; wr31<=w_6_703; wr32<=w_6_704; wr33<=w_6_705; wr34<=w_6_706; wr35<=w_6_707; wr36<=w_6_708; wr37<=w_6_709; wr38<=w_6_710; wr39<=w_6_711; wr40<=w_6_712; wr41<=w_6_713; wr42<=w_6_714; wr43<=w_6_715; wr44<=w_6_716; wr45<=w_6_717; wr46<=w_6_718; wr47<=w_6_719; wr48<=w_6_720; wr49<=w_6_721; wr50<=w_6_722; wr51<=w_6_723; wr52<=w_6_724; wr53<=w_6_725; wr54<=w_6_726; wr55<=w_6_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd104:
					begin
						wr0<=w_6_728; wr1<=w_6_729; wr2<=w_6_730; wr3<=w_6_731; wr4<=w_6_732; wr5<=w_6_733; wr6<=w_6_734; wr7<=w_6_735; wr8<=w_6_736; wr9<=w_6_737; wr10<=w_6_738; wr11<=w_6_739; wr12<=w_6_740; wr13<=w_6_741; wr14<=w_6_742; wr15<=w_6_743; wr16<=w_6_744; wr17<=w_6_745; wr18<=w_6_746; wr19<=w_6_747; wr20<=w_6_748; wr21<=w_6_749; wr22<=w_6_750; wr23<=w_6_751; wr24<=w_6_752; wr25<=w_6_753; wr26<=w_6_754; wr27<=w_6_755; wr28<=w_6_756; wr29<=w_6_757; wr30<=w_6_758; wr31<=w_6_759; wr32<=w_6_760; wr33<=w_6_761; wr34<=w_6_762; wr35<=w_6_763; wr36<=w_6_764; wr37<=w_6_765; wr38<=w_6_766; wr39<=w_6_767; wr40<=w_6_768; wr41<=w_6_769; wr42<=w_6_770; wr43<=w_6_771; wr44<=w_6_772; wr45<=w_6_773; wr46<=w_6_774; wr47<=w_6_775; wr48<=w_6_776; wr49<=w_6_777; wr50<=w_6_778; wr51<=w_6_779; wr52<=w_6_780; wr53<=w_6_781; wr54<=w_6_782; wr55<=w_6_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd105:
					begin
						bias_p<=px_784;
						bias_w<=w_6_784;
						select<=select+1;
					end
				8'd106:
					begin
						wr0<=w_7_0; wr1<=w_7_1; wr2<=w_7_2; wr3<=w_7_3; wr4<=w_7_4; wr5<=w_7_5; wr6<=w_7_6; wr7<=w_7_7; wr8<=w_7_8; wr9<=w_7_9; wr10<=w_7_10; wr11<=w_7_11; wr12<=w_7_12; wr13<=w_7_13; wr14<=w_7_14; wr15<=w_7_15; wr16<=w_7_16; wr17<=w_7_17; wr18<=w_7_18; wr19<=w_7_19; wr20<=w_7_20; wr21<=w_7_21; wr22<=w_7_22; wr23<=w_7_23; wr24<=w_7_24; wr25<=w_7_25; wr26<=w_7_26; wr27<=w_7_27; wr28<=w_7_28; wr29<=w_7_29; wr30<=w_7_30; wr31<=w_7_31; wr32<=w_7_32; wr33<=w_7_33; wr34<=w_7_34; wr35<=w_7_35; wr36<=w_7_36; wr37<=w_7_37; wr38<=w_7_38; wr39<=w_7_39; wr40<=w_7_40; wr41<=w_7_41; wr42<=w_7_42; wr43<=w_7_43; wr44<=w_7_44; wr45<=w_7_45; wr46<=w_7_46; wr47<=w_7_47; wr48<=w_7_48; wr49<=w_7_49; wr50<=w_7_50; wr51<=w_7_51; wr52<=w_7_52; wr53<=w_7_53; wr54<=w_7_54; wr55<=w_7_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd107:
					begin
						wr0<=w_7_56; wr1<=w_7_57; wr2<=w_7_58; wr3<=w_7_59; wr4<=w_7_60; wr5<=w_7_61; wr6<=w_7_62; wr7<=w_7_63; wr8<=w_7_64; wr9<=w_7_65; wr10<=w_7_66; wr11<=w_7_67; wr12<=w_7_68; wr13<=w_7_69; wr14<=w_7_70; wr15<=w_7_71; wr16<=w_7_72; wr17<=w_7_73; wr18<=w_7_74; wr19<=w_7_75; wr20<=w_7_76; wr21<=w_7_77; wr22<=w_7_78; wr23<=w_7_79; wr24<=w_7_80; wr25<=w_7_81; wr26<=w_7_82; wr27<=w_7_83; wr28<=w_7_84; wr29<=w_7_85; wr30<=w_7_86; wr31<=w_7_87; wr32<=w_7_88; wr33<=w_7_89; wr34<=w_7_90; wr35<=w_7_91; wr36<=w_7_92; wr37<=w_7_93; wr38<=w_7_94; wr39<=w_7_95; wr40<=w_7_96; wr41<=w_7_97; wr42<=w_7_98; wr43<=w_7_99; wr44<=w_7_100; wr45<=w_7_101; wr46<=w_7_102; wr47<=w_7_103; wr48<=w_7_104; wr49<=w_7_105; wr50<=w_7_106; wr51<=w_7_107; wr52<=w_7_108; wr53<=w_7_109; wr54<=w_7_110; wr55<=w_7_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd108:
					begin
						wr0<=w_7_112; wr1<=w_7_113; wr2<=w_7_114; wr3<=w_7_115; wr4<=w_7_116; wr5<=w_7_117; wr6<=w_7_118; wr7<=w_7_119; wr8<=w_7_120; wr9<=w_7_121; wr10<=w_7_122; wr11<=w_7_123; wr12<=w_7_124; wr13<=w_7_125; wr14<=w_7_126; wr15<=w_7_127; wr16<=w_7_128; wr17<=w_7_129; wr18<=w_7_130; wr19<=w_7_131; wr20<=w_7_132; wr21<=w_7_133; wr22<=w_7_134; wr23<=w_7_135; wr24<=w_7_136; wr25<=w_7_137; wr26<=w_7_138; wr27<=w_7_139; wr28<=w_7_140; wr29<=w_7_141; wr30<=w_7_142; wr31<=w_7_143; wr32<=w_7_144; wr33<=w_7_145; wr34<=w_7_146; wr35<=w_7_147; wr36<=w_7_148; wr37<=w_7_149; wr38<=w_7_150; wr39<=w_7_151; wr40<=w_7_152; wr41<=w_7_153; wr42<=w_7_154; wr43<=w_7_155; wr44<=w_7_156; wr45<=w_7_157; wr46<=w_7_158; wr47<=w_7_159; wr48<=w_7_160; wr49<=w_7_161; wr50<=w_7_162; wr51<=w_7_163; wr52<=w_7_164; wr53<=w_7_165; wr54<=w_7_166; wr55<=w_7_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd109:
					begin
						wr0<=w_7_168; wr1<=w_7_169; wr2<=w_7_170; wr3<=w_7_171; wr4<=w_7_172; wr5<=w_7_173; wr6<=w_7_174; wr7<=w_7_175; wr8<=w_7_176; wr9<=w_7_177; wr10<=w_7_178; wr11<=w_7_179; wr12<=w_7_180; wr13<=w_7_181; wr14<=w_7_182; wr15<=w_7_183; wr16<=w_7_184; wr17<=w_7_185; wr18<=w_7_186; wr19<=w_7_187; wr20<=w_7_188; wr21<=w_7_189; wr22<=w_7_190; wr23<=w_7_191; wr24<=w_7_192; wr25<=w_7_193; wr26<=w_7_194; wr27<=w_7_195; wr28<=w_7_196; wr29<=w_7_197; wr30<=w_7_198; wr31<=w_7_199; wr32<=w_7_200; wr33<=w_7_201; wr34<=w_7_202; wr35<=w_7_203; wr36<=w_7_204; wr37<=w_7_205; wr38<=w_7_206; wr39<=w_7_207; wr40<=w_7_208; wr41<=w_7_209; wr42<=w_7_210; wr43<=w_7_211; wr44<=w_7_212; wr45<=w_7_213; wr46<=w_7_214; wr47<=w_7_215; wr48<=w_7_216; wr49<=w_7_217; wr50<=w_7_218; wr51<=w_7_219; wr52<=w_7_220; wr53<=w_7_221; wr54<=w_7_222; wr55<=w_7_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd110:
					begin
						wr0<=w_7_224; wr1<=w_7_225; wr2<=w_7_226; wr3<=w_7_227; wr4<=w_7_228; wr5<=w_7_229; wr6<=w_7_230; wr7<=w_7_231; wr8<=w_7_232; wr9<=w_7_233; wr10<=w_7_234; wr11<=w_7_235; wr12<=w_7_236; wr13<=w_7_237; wr14<=w_7_238; wr15<=w_7_239; wr16<=w_7_240; wr17<=w_7_241; wr18<=w_7_242; wr19<=w_7_243; wr20<=w_7_244; wr21<=w_7_245; wr22<=w_7_246; wr23<=w_7_247; wr24<=w_7_248; wr25<=w_7_249; wr26<=w_7_250; wr27<=w_7_251; wr28<=w_7_252; wr29<=w_7_253; wr30<=w_7_254; wr31<=w_7_255; wr32<=w_7_256; wr33<=w_7_257; wr34<=w_7_258; wr35<=w_7_259; wr36<=w_7_260; wr37<=w_7_261; wr38<=w_7_262; wr39<=w_7_263; wr40<=w_7_264; wr41<=w_7_265; wr42<=w_7_266; wr43<=w_7_267; wr44<=w_7_268; wr45<=w_7_269; wr46<=w_7_270; wr47<=w_7_271; wr48<=w_7_272; wr49<=w_7_273; wr50<=w_7_274; wr51<=w_7_275; wr52<=w_7_276; wr53<=w_7_277; wr54<=w_7_278; wr55<=w_7_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd111:
					begin
						wr0<=w_7_280; wr1<=w_7_281; wr2<=w_7_282; wr3<=w_7_283; wr4<=w_7_284; wr5<=w_7_285; wr6<=w_7_286; wr7<=w_7_287; wr8<=w_7_288; wr9<=w_7_289; wr10<=w_7_290; wr11<=w_7_291; wr12<=w_7_292; wr13<=w_7_293; wr14<=w_7_294; wr15<=w_7_295; wr16<=w_7_296; wr17<=w_7_297; wr18<=w_7_298; wr19<=w_7_299; wr20<=w_7_300; wr21<=w_7_301; wr22<=w_7_302; wr23<=w_7_303; wr24<=w_7_304; wr25<=w_7_305; wr26<=w_7_306; wr27<=w_7_307; wr28<=w_7_308; wr29<=w_7_309; wr30<=w_7_310; wr31<=w_7_311; wr32<=w_7_312; wr33<=w_7_313; wr34<=w_7_314; wr35<=w_7_315; wr36<=w_7_316; wr37<=w_7_317; wr38<=w_7_318; wr39<=w_7_319; wr40<=w_7_320; wr41<=w_7_321; wr42<=w_7_322; wr43<=w_7_323; wr44<=w_7_324; wr45<=w_7_325; wr46<=w_7_326; wr47<=w_7_327; wr48<=w_7_328; wr49<=w_7_329; wr50<=w_7_330; wr51<=w_7_331; wr52<=w_7_332; wr53<=w_7_333; wr54<=w_7_334; wr55<=w_7_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd112:
					begin
						wr0<=w_7_336; wr1<=w_7_337; wr2<=w_7_338; wr3<=w_7_339; wr4<=w_7_340; wr5<=w_7_341; wr6<=w_7_342; wr7<=w_7_343; wr8<=w_7_344; wr9<=w_7_345; wr10<=w_7_346; wr11<=w_7_347; wr12<=w_7_348; wr13<=w_7_349; wr14<=w_7_350; wr15<=w_7_351; wr16<=w_7_352; wr17<=w_7_353; wr18<=w_7_354; wr19<=w_7_355; wr20<=w_7_356; wr21<=w_7_357; wr22<=w_7_358; wr23<=w_7_359; wr24<=w_7_360; wr25<=w_7_361; wr26<=w_7_362; wr27<=w_7_363; wr28<=w_7_364; wr29<=w_7_365; wr30<=w_7_366; wr31<=w_7_367; wr32<=w_7_368; wr33<=w_7_369; wr34<=w_7_370; wr35<=w_7_371; wr36<=w_7_372; wr37<=w_7_373; wr38<=w_7_374; wr39<=w_7_375; wr40<=w_7_376; wr41<=w_7_377; wr42<=w_7_378; wr43<=w_7_379; wr44<=w_7_380; wr45<=w_7_381; wr46<=w_7_382; wr47<=w_7_383; wr48<=w_7_384; wr49<=w_7_385; wr50<=w_7_386; wr51<=w_7_387; wr52<=w_7_388; wr53<=w_7_389; wr54<=w_7_390; wr55<=w_7_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd113:
					begin
						wr0<=w_7_392; wr1<=w_7_393; wr2<=w_7_394; wr3<=w_7_395; wr4<=w_7_396; wr5<=w_7_397; wr6<=w_7_398; wr7<=w_7_399; wr8<=w_7_400; wr9<=w_7_401; wr10<=w_7_402; wr11<=w_7_403; wr12<=w_7_404; wr13<=w_7_405; wr14<=w_7_406; wr15<=w_7_407; wr16<=w_7_408; wr17<=w_7_409; wr18<=w_7_410; wr19<=w_7_411; wr20<=w_7_412; wr21<=w_7_413; wr22<=w_7_414; wr23<=w_7_415; wr24<=w_7_416; wr25<=w_7_417; wr26<=w_7_418; wr27<=w_7_419; wr28<=w_7_420; wr29<=w_7_421; wr30<=w_7_422; wr31<=w_7_423; wr32<=w_7_424; wr33<=w_7_425; wr34<=w_7_426; wr35<=w_7_427; wr36<=w_7_428; wr37<=w_7_429; wr38<=w_7_430; wr39<=w_7_431; wr40<=w_7_432; wr41<=w_7_433; wr42<=w_7_434; wr43<=w_7_435; wr44<=w_7_436; wr45<=w_7_437; wr46<=w_7_438; wr47<=w_7_439; wr48<=w_7_440; wr49<=w_7_441; wr50<=w_7_442; wr51<=w_7_443; wr52<=w_7_444; wr53<=w_7_445; wr54<=w_7_446; wr55<=w_7_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd114:
					begin
						wr0<=w_7_448; wr1<=w_7_449; wr2<=w_7_450; wr3<=w_7_451; wr4<=w_7_452; wr5<=w_7_453; wr6<=w_7_454; wr7<=w_7_455; wr8<=w_7_456; wr9<=w_7_457; wr10<=w_7_458; wr11<=w_7_459; wr12<=w_7_460; wr13<=w_7_461; wr14<=w_7_462; wr15<=w_7_463; wr16<=w_7_464; wr17<=w_7_465; wr18<=w_7_466; wr19<=w_7_467; wr20<=w_7_468; wr21<=w_7_469; wr22<=w_7_470; wr23<=w_7_471; wr24<=w_7_472; wr25<=w_7_473; wr26<=w_7_474; wr27<=w_7_475; wr28<=w_7_476; wr29<=w_7_477; wr30<=w_7_478; wr31<=w_7_479; wr32<=w_7_480; wr33<=w_7_481; wr34<=w_7_482; wr35<=w_7_483; wr36<=w_7_484; wr37<=w_7_485; wr38<=w_7_486; wr39<=w_7_487; wr40<=w_7_488; wr41<=w_7_489; wr42<=w_7_490; wr43<=w_7_491; wr44<=w_7_492; wr45<=w_7_493; wr46<=w_7_494; wr47<=w_7_495; wr48<=w_7_496; wr49<=w_7_497; wr50<=w_7_498; wr51<=w_7_499; wr52<=w_7_500; wr53<=w_7_501; wr54<=w_7_502; wr55<=w_7_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd115:
					begin
						wr0<=w_7_504; wr1<=w_7_505; wr2<=w_7_506; wr3<=w_7_507; wr4<=w_7_508; wr5<=w_7_509; wr6<=w_7_510; wr7<=w_7_511; wr8<=w_7_512; wr9<=w_7_513; wr10<=w_7_514; wr11<=w_7_515; wr12<=w_7_516; wr13<=w_7_517; wr14<=w_7_518; wr15<=w_7_519; wr16<=w_7_520; wr17<=w_7_521; wr18<=w_7_522; wr19<=w_7_523; wr20<=w_7_524; wr21<=w_7_525; wr22<=w_7_526; wr23<=w_7_527; wr24<=w_7_528; wr25<=w_7_529; wr26<=w_7_530; wr27<=w_7_531; wr28<=w_7_532; wr29<=w_7_533; wr30<=w_7_534; wr31<=w_7_535; wr32<=w_7_536; wr33<=w_7_537; wr34<=w_7_538; wr35<=w_7_539; wr36<=w_7_540; wr37<=w_7_541; wr38<=w_7_542; wr39<=w_7_543; wr40<=w_7_544; wr41<=w_7_545; wr42<=w_7_546; wr43<=w_7_547; wr44<=w_7_548; wr45<=w_7_549; wr46<=w_7_550; wr47<=w_7_551; wr48<=w_7_552; wr49<=w_7_553; wr50<=w_7_554; wr51<=w_7_555; wr52<=w_7_556; wr53<=w_7_557; wr54<=w_7_558; wr55<=w_7_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd116:
					begin
						wr0<=w_7_560; wr1<=w_7_561; wr2<=w_7_562; wr3<=w_7_563; wr4<=w_7_564; wr5<=w_7_565; wr6<=w_7_566; wr7<=w_7_567; wr8<=w_7_568; wr9<=w_7_569; wr10<=w_7_570; wr11<=w_7_571; wr12<=w_7_572; wr13<=w_7_573; wr14<=w_7_574; wr15<=w_7_575; wr16<=w_7_576; wr17<=w_7_577; wr18<=w_7_578; wr19<=w_7_579; wr20<=w_7_580; wr21<=w_7_581; wr22<=w_7_582; wr23<=w_7_583; wr24<=w_7_584; wr25<=w_7_585; wr26<=w_7_586; wr27<=w_7_587; wr28<=w_7_588; wr29<=w_7_589; wr30<=w_7_590; wr31<=w_7_591; wr32<=w_7_592; wr33<=w_7_593; wr34<=w_7_594; wr35<=w_7_595; wr36<=w_7_596; wr37<=w_7_597; wr38<=w_7_598; wr39<=w_7_599; wr40<=w_7_600; wr41<=w_7_601; wr42<=w_7_602; wr43<=w_7_603; wr44<=w_7_604; wr45<=w_7_605; wr46<=w_7_606; wr47<=w_7_607; wr48<=w_7_608; wr49<=w_7_609; wr50<=w_7_610; wr51<=w_7_611; wr52<=w_7_612; wr53<=w_7_613; wr54<=w_7_614; wr55<=w_7_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd117:
					begin
						wr0<=w_7_616; wr1<=w_7_617; wr2<=w_7_618; wr3<=w_7_619; wr4<=w_7_620; wr5<=w_7_621; wr6<=w_7_622; wr7<=w_7_623; wr8<=w_7_624; wr9<=w_7_625; wr10<=w_7_626; wr11<=w_7_627; wr12<=w_7_628; wr13<=w_7_629; wr14<=w_7_630; wr15<=w_7_631; wr16<=w_7_632; wr17<=w_7_633; wr18<=w_7_634; wr19<=w_7_635; wr20<=w_7_636; wr21<=w_7_637; wr22<=w_7_638; wr23<=w_7_639; wr24<=w_7_640; wr25<=w_7_641; wr26<=w_7_642; wr27<=w_7_643; wr28<=w_7_644; wr29<=w_7_645; wr30<=w_7_646; wr31<=w_7_647; wr32<=w_7_648; wr33<=w_7_649; wr34<=w_7_650; wr35<=w_7_651; wr36<=w_7_652; wr37<=w_7_653; wr38<=w_7_654; wr39<=w_7_655; wr40<=w_7_656; wr41<=w_7_657; wr42<=w_7_658; wr43<=w_7_659; wr44<=w_7_660; wr45<=w_7_661; wr46<=w_7_662; wr47<=w_7_663; wr48<=w_7_664; wr49<=w_7_665; wr50<=w_7_666; wr51<=w_7_667; wr52<=w_7_668; wr53<=w_7_669; wr54<=w_7_670; wr55<=w_7_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd118:
					begin
						wr0<=w_7_672; wr1<=w_7_673; wr2<=w_7_674; wr3<=w_7_675; wr4<=w_7_676; wr5<=w_7_677; wr6<=w_7_678; wr7<=w_7_679; wr8<=w_7_680; wr9<=w_7_681; wr10<=w_7_682; wr11<=w_7_683; wr12<=w_7_684; wr13<=w_7_685; wr14<=w_7_686; wr15<=w_7_687; wr16<=w_7_688; wr17<=w_7_689; wr18<=w_7_690; wr19<=w_7_691; wr20<=w_7_692; wr21<=w_7_693; wr22<=w_7_694; wr23<=w_7_695; wr24<=w_7_696; wr25<=w_7_697; wr26<=w_7_698; wr27<=w_7_699; wr28<=w_7_700; wr29<=w_7_701; wr30<=w_7_702; wr31<=w_7_703; wr32<=w_7_704; wr33<=w_7_705; wr34<=w_7_706; wr35<=w_7_707; wr36<=w_7_708; wr37<=w_7_709; wr38<=w_7_710; wr39<=w_7_711; wr40<=w_7_712; wr41<=w_7_713; wr42<=w_7_714; wr43<=w_7_715; wr44<=w_7_716; wr45<=w_7_717; wr46<=w_7_718; wr47<=w_7_719; wr48<=w_7_720; wr49<=w_7_721; wr50<=w_7_722; wr51<=w_7_723; wr52<=w_7_724; wr53<=w_7_725; wr54<=w_7_726; wr55<=w_7_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd119:
					begin
						wr0<=w_7_728; wr1<=w_7_729; wr2<=w_7_730; wr3<=w_7_731; wr4<=w_7_732; wr5<=w_7_733; wr6<=w_7_734; wr7<=w_7_735; wr8<=w_7_736; wr9<=w_7_737; wr10<=w_7_738; wr11<=w_7_739; wr12<=w_7_740; wr13<=w_7_741; wr14<=w_7_742; wr15<=w_7_743; wr16<=w_7_744; wr17<=w_7_745; wr18<=w_7_746; wr19<=w_7_747; wr20<=w_7_748; wr21<=w_7_749; wr22<=w_7_750; wr23<=w_7_751; wr24<=w_7_752; wr25<=w_7_753; wr26<=w_7_754; wr27<=w_7_755; wr28<=w_7_756; wr29<=w_7_757; wr30<=w_7_758; wr31<=w_7_759; wr32<=w_7_760; wr33<=w_7_761; wr34<=w_7_762; wr35<=w_7_763; wr36<=w_7_764; wr37<=w_7_765; wr38<=w_7_766; wr39<=w_7_767; wr40<=w_7_768; wr41<=w_7_769; wr42<=w_7_770; wr43<=w_7_771; wr44<=w_7_772; wr45<=w_7_773; wr46<=w_7_774; wr47<=w_7_775; wr48<=w_7_776; wr49<=w_7_777; wr50<=w_7_778; wr51<=w_7_779; wr52<=w_7_780; wr53<=w_7_781; wr54<=w_7_782; wr55<=w_7_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd120:
					begin
						bias_p<=px_784;
						bias_w<=w_7_784;
						select<=select+1;
					end
				8'd121:
					begin
						wr0<=w_8_0; wr1<=w_8_1; wr2<=w_8_2; wr3<=w_8_3; wr4<=w_8_4; wr5<=w_8_5; wr6<=w_8_6; wr7<=w_8_7; wr8<=w_8_8; wr9<=w_8_9; wr10<=w_8_10; wr11<=w_8_11; wr12<=w_8_12; wr13<=w_8_13; wr14<=w_8_14; wr15<=w_8_15; wr16<=w_8_16; wr17<=w_8_17; wr18<=w_8_18; wr19<=w_8_19; wr20<=w_8_20; wr21<=w_8_21; wr22<=w_8_22; wr23<=w_8_23; wr24<=w_8_24; wr25<=w_8_25; wr26<=w_8_26; wr27<=w_8_27; wr28<=w_8_28; wr29<=w_8_29; wr30<=w_8_30; wr31<=w_8_31; wr32<=w_8_32; wr33<=w_8_33; wr34<=w_8_34; wr35<=w_8_35; wr36<=w_8_36; wr37<=w_8_37; wr38<=w_8_38; wr39<=w_8_39; wr40<=w_8_40; wr41<=w_8_41; wr42<=w_8_42; wr43<=w_8_43; wr44<=w_8_44; wr45<=w_8_45; wr46<=w_8_46; wr47<=w_8_47; wr48<=w_8_48; wr49<=w_8_49; wr50<=w_8_50; wr51<=w_8_51; wr52<=w_8_52; wr53<=w_8_53; wr54<=w_8_54; wr55<=w_8_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd122:
					begin
						wr0<=w_8_56; wr1<=w_8_57; wr2<=w_8_58; wr3<=w_8_59; wr4<=w_8_60; wr5<=w_8_61; wr6<=w_8_62; wr7<=w_8_63; wr8<=w_8_64; wr9<=w_8_65; wr10<=w_8_66; wr11<=w_8_67; wr12<=w_8_68; wr13<=w_8_69; wr14<=w_8_70; wr15<=w_8_71; wr16<=w_8_72; wr17<=w_8_73; wr18<=w_8_74; wr19<=w_8_75; wr20<=w_8_76; wr21<=w_8_77; wr22<=w_8_78; wr23<=w_8_79; wr24<=w_8_80; wr25<=w_8_81; wr26<=w_8_82; wr27<=w_8_83; wr28<=w_8_84; wr29<=w_8_85; wr30<=w_8_86; wr31<=w_8_87; wr32<=w_8_88; wr33<=w_8_89; wr34<=w_8_90; wr35<=w_8_91; wr36<=w_8_92; wr37<=w_8_93; wr38<=w_8_94; wr39<=w_8_95; wr40<=w_8_96; wr41<=w_8_97; wr42<=w_8_98; wr43<=w_8_99; wr44<=w_8_100; wr45<=w_8_101; wr46<=w_8_102; wr47<=w_8_103; wr48<=w_8_104; wr49<=w_8_105; wr50<=w_8_106; wr51<=w_8_107; wr52<=w_8_108; wr53<=w_8_109; wr54<=w_8_110; wr55<=w_8_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd123:
					begin
						wr0<=w_8_112; wr1<=w_8_113; wr2<=w_8_114; wr3<=w_8_115; wr4<=w_8_116; wr5<=w_8_117; wr6<=w_8_118; wr7<=w_8_119; wr8<=w_8_120; wr9<=w_8_121; wr10<=w_8_122; wr11<=w_8_123; wr12<=w_8_124; wr13<=w_8_125; wr14<=w_8_126; wr15<=w_8_127; wr16<=w_8_128; wr17<=w_8_129; wr18<=w_8_130; wr19<=w_8_131; wr20<=w_8_132; wr21<=w_8_133; wr22<=w_8_134; wr23<=w_8_135; wr24<=w_8_136; wr25<=w_8_137; wr26<=w_8_138; wr27<=w_8_139; wr28<=w_8_140; wr29<=w_8_141; wr30<=w_8_142; wr31<=w_8_143; wr32<=w_8_144; wr33<=w_8_145; wr34<=w_8_146; wr35<=w_8_147; wr36<=w_8_148; wr37<=w_8_149; wr38<=w_8_150; wr39<=w_8_151; wr40<=w_8_152; wr41<=w_8_153; wr42<=w_8_154; wr43<=w_8_155; wr44<=w_8_156; wr45<=w_8_157; wr46<=w_8_158; wr47<=w_8_159; wr48<=w_8_160; wr49<=w_8_161; wr50<=w_8_162; wr51<=w_8_163; wr52<=w_8_164; wr53<=w_8_165; wr54<=w_8_166; wr55<=w_8_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd124:
					begin
						wr0<=w_8_168; wr1<=w_8_169; wr2<=w_8_170; wr3<=w_8_171; wr4<=w_8_172; wr5<=w_8_173; wr6<=w_8_174; wr7<=w_8_175; wr8<=w_8_176; wr9<=w_8_177; wr10<=w_8_178; wr11<=w_8_179; wr12<=w_8_180; wr13<=w_8_181; wr14<=w_8_182; wr15<=w_8_183; wr16<=w_8_184; wr17<=w_8_185; wr18<=w_8_186; wr19<=w_8_187; wr20<=w_8_188; wr21<=w_8_189; wr22<=w_8_190; wr23<=w_8_191; wr24<=w_8_192; wr25<=w_8_193; wr26<=w_8_194; wr27<=w_8_195; wr28<=w_8_196; wr29<=w_8_197; wr30<=w_8_198; wr31<=w_8_199; wr32<=w_8_200; wr33<=w_8_201; wr34<=w_8_202; wr35<=w_8_203; wr36<=w_8_204; wr37<=w_8_205; wr38<=w_8_206; wr39<=w_8_207; wr40<=w_8_208; wr41<=w_8_209; wr42<=w_8_210; wr43<=w_8_211; wr44<=w_8_212; wr45<=w_8_213; wr46<=w_8_214; wr47<=w_8_215; wr48<=w_8_216; wr49<=w_8_217; wr50<=w_8_218; wr51<=w_8_219; wr52<=w_8_220; wr53<=w_8_221; wr54<=w_8_222; wr55<=w_8_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd125:
					begin
						wr0<=w_8_224; wr1<=w_8_225; wr2<=w_8_226; wr3<=w_8_227; wr4<=w_8_228; wr5<=w_8_229; wr6<=w_8_230; wr7<=w_8_231; wr8<=w_8_232; wr9<=w_8_233; wr10<=w_8_234; wr11<=w_8_235; wr12<=w_8_236; wr13<=w_8_237; wr14<=w_8_238; wr15<=w_8_239; wr16<=w_8_240; wr17<=w_8_241; wr18<=w_8_242; wr19<=w_8_243; wr20<=w_8_244; wr21<=w_8_245; wr22<=w_8_246; wr23<=w_8_247; wr24<=w_8_248; wr25<=w_8_249; wr26<=w_8_250; wr27<=w_8_251; wr28<=w_8_252; wr29<=w_8_253; wr30<=w_8_254; wr31<=w_8_255; wr32<=w_8_256; wr33<=w_8_257; wr34<=w_8_258; wr35<=w_8_259; wr36<=w_8_260; wr37<=w_8_261; wr38<=w_8_262; wr39<=w_8_263; wr40<=w_8_264; wr41<=w_8_265; wr42<=w_8_266; wr43<=w_8_267; wr44<=w_8_268; wr45<=w_8_269; wr46<=w_8_270; wr47<=w_8_271; wr48<=w_8_272; wr49<=w_8_273; wr50<=w_8_274; wr51<=w_8_275; wr52<=w_8_276; wr53<=w_8_277; wr54<=w_8_278; wr55<=w_8_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd126:
					begin
						wr0<=w_8_280; wr1<=w_8_281; wr2<=w_8_282; wr3<=w_8_283; wr4<=w_8_284; wr5<=w_8_285; wr6<=w_8_286; wr7<=w_8_287; wr8<=w_8_288; wr9<=w_8_289; wr10<=w_8_290; wr11<=w_8_291; wr12<=w_8_292; wr13<=w_8_293; wr14<=w_8_294; wr15<=w_8_295; wr16<=w_8_296; wr17<=w_8_297; wr18<=w_8_298; wr19<=w_8_299; wr20<=w_8_300; wr21<=w_8_301; wr22<=w_8_302; wr23<=w_8_303; wr24<=w_8_304; wr25<=w_8_305; wr26<=w_8_306; wr27<=w_8_307; wr28<=w_8_308; wr29<=w_8_309; wr30<=w_8_310; wr31<=w_8_311; wr32<=w_8_312; wr33<=w_8_313; wr34<=w_8_314; wr35<=w_8_315; wr36<=w_8_316; wr37<=w_8_317; wr38<=w_8_318; wr39<=w_8_319; wr40<=w_8_320; wr41<=w_8_321; wr42<=w_8_322; wr43<=w_8_323; wr44<=w_8_324; wr45<=w_8_325; wr46<=w_8_326; wr47<=w_8_327; wr48<=w_8_328; wr49<=w_8_329; wr50<=w_8_330; wr51<=w_8_331; wr52<=w_8_332; wr53<=w_8_333; wr54<=w_8_334; wr55<=w_8_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd127:
					begin
						wr0<=w_8_336; wr1<=w_8_337; wr2<=w_8_338; wr3<=w_8_339; wr4<=w_8_340; wr5<=w_8_341; wr6<=w_8_342; wr7<=w_8_343; wr8<=w_8_344; wr9<=w_8_345; wr10<=w_8_346; wr11<=w_8_347; wr12<=w_8_348; wr13<=w_8_349; wr14<=w_8_350; wr15<=w_8_351; wr16<=w_8_352; wr17<=w_8_353; wr18<=w_8_354; wr19<=w_8_355; wr20<=w_8_356; wr21<=w_8_357; wr22<=w_8_358; wr23<=w_8_359; wr24<=w_8_360; wr25<=w_8_361; wr26<=w_8_362; wr27<=w_8_363; wr28<=w_8_364; wr29<=w_8_365; wr30<=w_8_366; wr31<=w_8_367; wr32<=w_8_368; wr33<=w_8_369; wr34<=w_8_370; wr35<=w_8_371; wr36<=w_8_372; wr37<=w_8_373; wr38<=w_8_374; wr39<=w_8_375; wr40<=w_8_376; wr41<=w_8_377; wr42<=w_8_378; wr43<=w_8_379; wr44<=w_8_380; wr45<=w_8_381; wr46<=w_8_382; wr47<=w_8_383; wr48<=w_8_384; wr49<=w_8_385; wr50<=w_8_386; wr51<=w_8_387; wr52<=w_8_388; wr53<=w_8_389; wr54<=w_8_390; wr55<=w_8_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd128:
					begin
						wr0<=w_8_392; wr1<=w_8_393; wr2<=w_8_394; wr3<=w_8_395; wr4<=w_8_396; wr5<=w_8_397; wr6<=w_8_398; wr7<=w_8_399; wr8<=w_8_400; wr9<=w_8_401; wr10<=w_8_402; wr11<=w_8_403; wr12<=w_8_404; wr13<=w_8_405; wr14<=w_8_406; wr15<=w_8_407; wr16<=w_8_408; wr17<=w_8_409; wr18<=w_8_410; wr19<=w_8_411; wr20<=w_8_412; wr21<=w_8_413; wr22<=w_8_414; wr23<=w_8_415; wr24<=w_8_416; wr25<=w_8_417; wr26<=w_8_418; wr27<=w_8_419; wr28<=w_8_420; wr29<=w_8_421; wr30<=w_8_422; wr31<=w_8_423; wr32<=w_8_424; wr33<=w_8_425; wr34<=w_8_426; wr35<=w_8_427; wr36<=w_8_428; wr37<=w_8_429; wr38<=w_8_430; wr39<=w_8_431; wr40<=w_8_432; wr41<=w_8_433; wr42<=w_8_434; wr43<=w_8_435; wr44<=w_8_436; wr45<=w_8_437; wr46<=w_8_438; wr47<=w_8_439; wr48<=w_8_440; wr49<=w_8_441; wr50<=w_8_442; wr51<=w_8_443; wr52<=w_8_444; wr53<=w_8_445; wr54<=w_8_446; wr55<=w_8_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd129:
					begin
						wr0<=w_8_448; wr1<=w_8_449; wr2<=w_8_450; wr3<=w_8_451; wr4<=w_8_452; wr5<=w_8_453; wr6<=w_8_454; wr7<=w_8_455; wr8<=w_8_456; wr9<=w_8_457; wr10<=w_8_458; wr11<=w_8_459; wr12<=w_8_460; wr13<=w_8_461; wr14<=w_8_462; wr15<=w_8_463; wr16<=w_8_464; wr17<=w_8_465; wr18<=w_8_466; wr19<=w_8_467; wr20<=w_8_468; wr21<=w_8_469; wr22<=w_8_470; wr23<=w_8_471; wr24<=w_8_472; wr25<=w_8_473; wr26<=w_8_474; wr27<=w_8_475; wr28<=w_8_476; wr29<=w_8_477; wr30<=w_8_478; wr31<=w_8_479; wr32<=w_8_480; wr33<=w_8_481; wr34<=w_8_482; wr35<=w_8_483; wr36<=w_8_484; wr37<=w_8_485; wr38<=w_8_486; wr39<=w_8_487; wr40<=w_8_488; wr41<=w_8_489; wr42<=w_8_490; wr43<=w_8_491; wr44<=w_8_492; wr45<=w_8_493; wr46<=w_8_494; wr47<=w_8_495; wr48<=w_8_496; wr49<=w_8_497; wr50<=w_8_498; wr51<=w_8_499; wr52<=w_8_500; wr53<=w_8_501; wr54<=w_8_502; wr55<=w_8_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd130:
					begin
						wr0<=w_8_504; wr1<=w_8_505; wr2<=w_8_506; wr3<=w_8_507; wr4<=w_8_508; wr5<=w_8_509; wr6<=w_8_510; wr7<=w_8_511; wr8<=w_8_512; wr9<=w_8_513; wr10<=w_8_514; wr11<=w_8_515; wr12<=w_8_516; wr13<=w_8_517; wr14<=w_8_518; wr15<=w_8_519; wr16<=w_8_520; wr17<=w_8_521; wr18<=w_8_522; wr19<=w_8_523; wr20<=w_8_524; wr21<=w_8_525; wr22<=w_8_526; wr23<=w_8_527; wr24<=w_8_528; wr25<=w_8_529; wr26<=w_8_530; wr27<=w_8_531; wr28<=w_8_532; wr29<=w_8_533; wr30<=w_8_534; wr31<=w_8_535; wr32<=w_8_536; wr33<=w_8_537; wr34<=w_8_538; wr35<=w_8_539; wr36<=w_8_540; wr37<=w_8_541; wr38<=w_8_542; wr39<=w_8_543; wr40<=w_8_544; wr41<=w_8_545; wr42<=w_8_546; wr43<=w_8_547; wr44<=w_8_548; wr45<=w_8_549; wr46<=w_8_550; wr47<=w_8_551; wr48<=w_8_552; wr49<=w_8_553; wr50<=w_8_554; wr51<=w_8_555; wr52<=w_8_556; wr53<=w_8_557; wr54<=w_8_558; wr55<=w_8_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd131:
					begin
						wr0<=w_8_560; wr1<=w_8_561; wr2<=w_8_562; wr3<=w_8_563; wr4<=w_8_564; wr5<=w_8_565; wr6<=w_8_566; wr7<=w_8_567; wr8<=w_8_568; wr9<=w_8_569; wr10<=w_8_570; wr11<=w_8_571; wr12<=w_8_572; wr13<=w_8_573; wr14<=w_8_574; wr15<=w_8_575; wr16<=w_8_576; wr17<=w_8_577; wr18<=w_8_578; wr19<=w_8_579; wr20<=w_8_580; wr21<=w_8_581; wr22<=w_8_582; wr23<=w_8_583; wr24<=w_8_584; wr25<=w_8_585; wr26<=w_8_586; wr27<=w_8_587; wr28<=w_8_588; wr29<=w_8_589; wr30<=w_8_590; wr31<=w_8_591; wr32<=w_8_592; wr33<=w_8_593; wr34<=w_8_594; wr35<=w_8_595; wr36<=w_8_596; wr37<=w_8_597; wr38<=w_8_598; wr39<=w_8_599; wr40<=w_8_600; wr41<=w_8_601; wr42<=w_8_602; wr43<=w_8_603; wr44<=w_8_604; wr45<=w_8_605; wr46<=w_8_606; wr47<=w_8_607; wr48<=w_8_608; wr49<=w_8_609; wr50<=w_8_610; wr51<=w_8_611; wr52<=w_8_612; wr53<=w_8_613; wr54<=w_8_614; wr55<=w_8_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd132:
					begin
						wr0<=w_8_616; wr1<=w_8_617; wr2<=w_8_618; wr3<=w_8_619; wr4<=w_8_620; wr5<=w_8_621; wr6<=w_8_622; wr7<=w_8_623; wr8<=w_8_624; wr9<=w_8_625; wr10<=w_8_626; wr11<=w_8_627; wr12<=w_8_628; wr13<=w_8_629; wr14<=w_8_630; wr15<=w_8_631; wr16<=w_8_632; wr17<=w_8_633; wr18<=w_8_634; wr19<=w_8_635; wr20<=w_8_636; wr21<=w_8_637; wr22<=w_8_638; wr23<=w_8_639; wr24<=w_8_640; wr25<=w_8_641; wr26<=w_8_642; wr27<=w_8_643; wr28<=w_8_644; wr29<=w_8_645; wr30<=w_8_646; wr31<=w_8_647; wr32<=w_8_648; wr33<=w_8_649; wr34<=w_8_650; wr35<=w_8_651; wr36<=w_8_652; wr37<=w_8_653; wr38<=w_8_654; wr39<=w_8_655; wr40<=w_8_656; wr41<=w_8_657; wr42<=w_8_658; wr43<=w_8_659; wr44<=w_8_660; wr45<=w_8_661; wr46<=w_8_662; wr47<=w_8_663; wr48<=w_8_664; wr49<=w_8_665; wr50<=w_8_666; wr51<=w_8_667; wr52<=w_8_668; wr53<=w_8_669; wr54<=w_8_670; wr55<=w_8_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd133:
					begin
						wr0<=w_8_672; wr1<=w_8_673; wr2<=w_8_674; wr3<=w_8_675; wr4<=w_8_676; wr5<=w_8_677; wr6<=w_8_678; wr7<=w_8_679; wr8<=w_8_680; wr9<=w_8_681; wr10<=w_8_682; wr11<=w_8_683; wr12<=w_8_684; wr13<=w_8_685; wr14<=w_8_686; wr15<=w_8_687; wr16<=w_8_688; wr17<=w_8_689; wr18<=w_8_690; wr19<=w_8_691; wr20<=w_8_692; wr21<=w_8_693; wr22<=w_8_694; wr23<=w_8_695; wr24<=w_8_696; wr25<=w_8_697; wr26<=w_8_698; wr27<=w_8_699; wr28<=w_8_700; wr29<=w_8_701; wr30<=w_8_702; wr31<=w_8_703; wr32<=w_8_704; wr33<=w_8_705; wr34<=w_8_706; wr35<=w_8_707; wr36<=w_8_708; wr37<=w_8_709; wr38<=w_8_710; wr39<=w_8_711; wr40<=w_8_712; wr41<=w_8_713; wr42<=w_8_714; wr43<=w_8_715; wr44<=w_8_716; wr45<=w_8_717; wr46<=w_8_718; wr47<=w_8_719; wr48<=w_8_720; wr49<=w_8_721; wr50<=w_8_722; wr51<=w_8_723; wr52<=w_8_724; wr53<=w_8_725; wr54<=w_8_726; wr55<=w_8_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd134:
					begin
						wr0<=w_8_728; wr1<=w_8_729; wr2<=w_8_730; wr3<=w_8_731; wr4<=w_8_732; wr5<=w_8_733; wr6<=w_8_734; wr7<=w_8_735; wr8<=w_8_736; wr9<=w_8_737; wr10<=w_8_738; wr11<=w_8_739; wr12<=w_8_740; wr13<=w_8_741; wr14<=w_8_742; wr15<=w_8_743; wr16<=w_8_744; wr17<=w_8_745; wr18<=w_8_746; wr19<=w_8_747; wr20<=w_8_748; wr21<=w_8_749; wr22<=w_8_750; wr23<=w_8_751; wr24<=w_8_752; wr25<=w_8_753; wr26<=w_8_754; wr27<=w_8_755; wr28<=w_8_756; wr29<=w_8_757; wr30<=w_8_758; wr31<=w_8_759; wr32<=w_8_760; wr33<=w_8_761; wr34<=w_8_762; wr35<=w_8_763; wr36<=w_8_764; wr37<=w_8_765; wr38<=w_8_766; wr39<=w_8_767; wr40<=w_8_768; wr41<=w_8_769; wr42<=w_8_770; wr43<=w_8_771; wr44<=w_8_772; wr45<=w_8_773; wr46<=w_8_774; wr47<=w_8_775; wr48<=w_8_776; wr49<=w_8_777; wr50<=w_8_778; wr51<=w_8_779; wr52<=w_8_780; wr53<=w_8_781; wr54<=w_8_782; wr55<=w_8_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd135:
					begin
						bias_p<=px_784;
						bias_w<=w_8_784;
						select<=select+1;
					end
				8'd136:
					begin
						wr0<=w_9_0; wr1<=w_9_1; wr2<=w_9_2; wr3<=w_9_3; wr4<=w_9_4; wr5<=w_9_5; wr6<=w_9_6; wr7<=w_9_7; wr8<=w_9_8; wr9<=w_9_9; wr10<=w_9_10; wr11<=w_9_11; wr12<=w_9_12; wr13<=w_9_13; wr14<=w_9_14; wr15<=w_9_15; wr16<=w_9_16; wr17<=w_9_17; wr18<=w_9_18; wr19<=w_9_19; wr20<=w_9_20; wr21<=w_9_21; wr22<=w_9_22; wr23<=w_9_23; wr24<=w_9_24; wr25<=w_9_25; wr26<=w_9_26; wr27<=w_9_27; wr28<=w_9_28; wr29<=w_9_29; wr30<=w_9_30; wr31<=w_9_31; wr32<=w_9_32; wr33<=w_9_33; wr34<=w_9_34; wr35<=w_9_35; wr36<=w_9_36; wr37<=w_9_37; wr38<=w_9_38; wr39<=w_9_39; wr40<=w_9_40; wr41<=w_9_41; wr42<=w_9_42; wr43<=w_9_43; wr44<=w_9_44; wr45<=w_9_45; wr46<=w_9_46; wr47<=w_9_47; wr48<=w_9_48; wr49<=w_9_49; wr50<=w_9_50; wr51<=w_9_51; wr52<=w_9_52; wr53<=w_9_53; wr54<=w_9_54; wr55<=w_9_55; 
						r0<=Pix_0; r1<=Pix_1; r2<=Pix_2; r3<=Pix_3; r4<=Pix_4; r5<=Pix_5; r6<=Pix_6; r7<=Pix_7; r8<=Pix_8; r9<=Pix_9; r10<=Pix_10; r11<=Pix_11; r12<=Pix_12; r13<=Pix_13; r14<=Pix_14; r15<=Pix_15; r16<=Pix_16; r17<=Pix_17; r18<=Pix_18; r19<=Pix_19; r20<=Pix_20; r21<=Pix_21; r22<=Pix_22; r23<=Pix_23; r24<=Pix_24; r25<=Pix_25; r26<=Pix_26; r27<=Pix_27; r28<=Pix_28; r29<=Pix_29; r30<=Pix_30; r31<=Pix_31; r32<=Pix_32; r33<=Pix_33; r34<=Pix_34; r35<=Pix_35; r36<=Pix_36; r37<=Pix_37; r38<=Pix_38; r39<=Pix_39; r40<=Pix_40; r41<=Pix_41; r42<=Pix_42; r43<=Pix_43; r44<=Pix_44; r45<=Pix_45; r46<=Pix_46; r47<=Pix_47; r48<=Pix_48; r49<=Pix_49; r50<=Pix_50; r51<=Pix_51; r52<=Pix_52; r53<=Pix_53; r54<=Pix_54; r55<=Pix_55; 
						select<=select+1;
					end
				8'd137:
					begin
						wr0<=w_9_56; wr1<=w_9_57; wr2<=w_9_58; wr3<=w_9_59; wr4<=w_9_60; wr5<=w_9_61; wr6<=w_9_62; wr7<=w_9_63; wr8<=w_9_64; wr9<=w_9_65; wr10<=w_9_66; wr11<=w_9_67; wr12<=w_9_68; wr13<=w_9_69; wr14<=w_9_70; wr15<=w_9_71; wr16<=w_9_72; wr17<=w_9_73; wr18<=w_9_74; wr19<=w_9_75; wr20<=w_9_76; wr21<=w_9_77; wr22<=w_9_78; wr23<=w_9_79; wr24<=w_9_80; wr25<=w_9_81; wr26<=w_9_82; wr27<=w_9_83; wr28<=w_9_84; wr29<=w_9_85; wr30<=w_9_86; wr31<=w_9_87; wr32<=w_9_88; wr33<=w_9_89; wr34<=w_9_90; wr35<=w_9_91; wr36<=w_9_92; wr37<=w_9_93; wr38<=w_9_94; wr39<=w_9_95; wr40<=w_9_96; wr41<=w_9_97; wr42<=w_9_98; wr43<=w_9_99; wr44<=w_9_100; wr45<=w_9_101; wr46<=w_9_102; wr47<=w_9_103; wr48<=w_9_104; wr49<=w_9_105; wr50<=w_9_106; wr51<=w_9_107; wr52<=w_9_108; wr53<=w_9_109; wr54<=w_9_110; wr55<=w_9_111; 
						r0<=Pix_56; r1<=Pix_57; r2<=Pix_58; r3<=Pix_59; r4<=Pix_60; r5<=Pix_61; r6<=Pix_62; r7<=Pix_63; r8<=Pix_64; r9<=Pix_65; r10<=Pix_66; r11<=Pix_67; r12<=Pix_68; r13<=Pix_69; r14<=Pix_70; r15<=Pix_71; r16<=Pix_72; r17<=Pix_73; r18<=Pix_74; r19<=Pix_75; r20<=Pix_76; r21<=Pix_77; r22<=Pix_78; r23<=Pix_79; r24<=Pix_80; r25<=Pix_81; r26<=Pix_82; r27<=Pix_83; r28<=Pix_84; r29<=Pix_85; r30<=Pix_86; r31<=Pix_87; r32<=Pix_88; r33<=Pix_89; r34<=Pix_90; r35<=Pix_91; r36<=Pix_92; r37<=Pix_93; r38<=Pix_94; r39<=Pix_95; r40<=Pix_96; r41<=Pix_97; r42<=Pix_98; r43<=Pix_99; r44<=Pix_100; r45<=Pix_101; r46<=Pix_102; r47<=Pix_103; r48<=Pix_104; r49<=Pix_105; r50<=Pix_106; r51<=Pix_107; r52<=Pix_108; r53<=Pix_109; r54<=Pix_110; r55<=Pix_111; 
						select<=select+1;
					end
				8'd138:
					begin
						wr0<=w_9_112; wr1<=w_9_113; wr2<=w_9_114; wr3<=w_9_115; wr4<=w_9_116; wr5<=w_9_117; wr6<=w_9_118; wr7<=w_9_119; wr8<=w_9_120; wr9<=w_9_121; wr10<=w_9_122; wr11<=w_9_123; wr12<=w_9_124; wr13<=w_9_125; wr14<=w_9_126; wr15<=w_9_127; wr16<=w_9_128; wr17<=w_9_129; wr18<=w_9_130; wr19<=w_9_131; wr20<=w_9_132; wr21<=w_9_133; wr22<=w_9_134; wr23<=w_9_135; wr24<=w_9_136; wr25<=w_9_137; wr26<=w_9_138; wr27<=w_9_139; wr28<=w_9_140; wr29<=w_9_141; wr30<=w_9_142; wr31<=w_9_143; wr32<=w_9_144; wr33<=w_9_145; wr34<=w_9_146; wr35<=w_9_147; wr36<=w_9_148; wr37<=w_9_149; wr38<=w_9_150; wr39<=w_9_151; wr40<=w_9_152; wr41<=w_9_153; wr42<=w_9_154; wr43<=w_9_155; wr44<=w_9_156; wr45<=w_9_157; wr46<=w_9_158; wr47<=w_9_159; wr48<=w_9_160; wr49<=w_9_161; wr50<=w_9_162; wr51<=w_9_163; wr52<=w_9_164; wr53<=w_9_165; wr54<=w_9_166; wr55<=w_9_167; 
						r0<=Pix_112; r1<=Pix_113; r2<=Pix_114; r3<=Pix_115; r4<=Pix_116; r5<=Pix_117; r6<=Pix_118; r7<=Pix_119; r8<=Pix_120; r9<=Pix_121; r10<=Pix_122; r11<=Pix_123; r12<=Pix_124; r13<=Pix_125; r14<=Pix_126; r15<=Pix_127; r16<=Pix_128; r17<=Pix_129; r18<=Pix_130; r19<=Pix_131; r20<=Pix_132; r21<=Pix_133; r22<=Pix_134; r23<=Pix_135; r24<=Pix_136; r25<=Pix_137; r26<=Pix_138; r27<=Pix_139; r28<=Pix_140; r29<=Pix_141; r30<=Pix_142; r31<=Pix_143; r32<=Pix_144; r33<=Pix_145; r34<=Pix_146; r35<=Pix_147; r36<=Pix_148; r37<=Pix_149; r38<=Pix_150; r39<=Pix_151; r40<=Pix_152; r41<=Pix_153; r42<=Pix_154; r43<=Pix_155; r44<=Pix_156; r45<=Pix_157; r46<=Pix_158; r47<=Pix_159; r48<=Pix_160; r49<=Pix_161; r50<=Pix_162; r51<=Pix_163; r52<=Pix_164; r53<=Pix_165; r54<=Pix_166; r55<=Pix_167; 
						select<=select+1;
					end
				8'd139:
					begin
						wr0<=w_9_168; wr1<=w_9_169; wr2<=w_9_170; wr3<=w_9_171; wr4<=w_9_172; wr5<=w_9_173; wr6<=w_9_174; wr7<=w_9_175; wr8<=w_9_176; wr9<=w_9_177; wr10<=w_9_178; wr11<=w_9_179; wr12<=w_9_180; wr13<=w_9_181; wr14<=w_9_182; wr15<=w_9_183; wr16<=w_9_184; wr17<=w_9_185; wr18<=w_9_186; wr19<=w_9_187; wr20<=w_9_188; wr21<=w_9_189; wr22<=w_9_190; wr23<=w_9_191; wr24<=w_9_192; wr25<=w_9_193; wr26<=w_9_194; wr27<=w_9_195; wr28<=w_9_196; wr29<=w_9_197; wr30<=w_9_198; wr31<=w_9_199; wr32<=w_9_200; wr33<=w_9_201; wr34<=w_9_202; wr35<=w_9_203; wr36<=w_9_204; wr37<=w_9_205; wr38<=w_9_206; wr39<=w_9_207; wr40<=w_9_208; wr41<=w_9_209; wr42<=w_9_210; wr43<=w_9_211; wr44<=w_9_212; wr45<=w_9_213; wr46<=w_9_214; wr47<=w_9_215; wr48<=w_9_216; wr49<=w_9_217; wr50<=w_9_218; wr51<=w_9_219; wr52<=w_9_220; wr53<=w_9_221; wr54<=w_9_222; wr55<=w_9_223; 
						r0<=Pix_168; r1<=Pix_169; r2<=Pix_170; r3<=Pix_171; r4<=Pix_172; r5<=Pix_173; r6<=Pix_174; r7<=Pix_175; r8<=Pix_176; r9<=Pix_177; r10<=Pix_178; r11<=Pix_179; r12<=Pix_180; r13<=Pix_181; r14<=Pix_182; r15<=Pix_183; r16<=Pix_184; r17<=Pix_185; r18<=Pix_186; r19<=Pix_187; r20<=Pix_188; r21<=Pix_189; r22<=Pix_190; r23<=Pix_191; r24<=Pix_192; r25<=Pix_193; r26<=Pix_194; r27<=Pix_195; r28<=Pix_196; r29<=Pix_197; r30<=Pix_198; r31<=Pix_199; r32<=Pix_200; r33<=Pix_201; r34<=Pix_202; r35<=Pix_203; r36<=Pix_204; r37<=Pix_205; r38<=Pix_206; r39<=Pix_207; r40<=Pix_208; r41<=Pix_209; r42<=Pix_210; r43<=Pix_211; r44<=Pix_212; r45<=Pix_213; r46<=Pix_214; r47<=Pix_215; r48<=Pix_216; r49<=Pix_217; r50<=Pix_218; r51<=Pix_219; r52<=Pix_220; r53<=Pix_221; r54<=Pix_222; r55<=Pix_223; 
						select<=select+1;
					end
				8'd140:
					begin
						wr0<=w_9_224; wr1<=w_9_225; wr2<=w_9_226; wr3<=w_9_227; wr4<=w_9_228; wr5<=w_9_229; wr6<=w_9_230; wr7<=w_9_231; wr8<=w_9_232; wr9<=w_9_233; wr10<=w_9_234; wr11<=w_9_235; wr12<=w_9_236; wr13<=w_9_237; wr14<=w_9_238; wr15<=w_9_239; wr16<=w_9_240; wr17<=w_9_241; wr18<=w_9_242; wr19<=w_9_243; wr20<=w_9_244; wr21<=w_9_245; wr22<=w_9_246; wr23<=w_9_247; wr24<=w_9_248; wr25<=w_9_249; wr26<=w_9_250; wr27<=w_9_251; wr28<=w_9_252; wr29<=w_9_253; wr30<=w_9_254; wr31<=w_9_255; wr32<=w_9_256; wr33<=w_9_257; wr34<=w_9_258; wr35<=w_9_259; wr36<=w_9_260; wr37<=w_9_261; wr38<=w_9_262; wr39<=w_9_263; wr40<=w_9_264; wr41<=w_9_265; wr42<=w_9_266; wr43<=w_9_267; wr44<=w_9_268; wr45<=w_9_269; wr46<=w_9_270; wr47<=w_9_271; wr48<=w_9_272; wr49<=w_9_273; wr50<=w_9_274; wr51<=w_9_275; wr52<=w_9_276; wr53<=w_9_277; wr54<=w_9_278; wr55<=w_9_279; 
						r0<=Pix_224; r1<=Pix_225; r2<=Pix_226; r3<=Pix_227; r4<=Pix_228; r5<=Pix_229; r6<=Pix_230; r7<=Pix_231; r8<=Pix_232; r9<=Pix_233; r10<=Pix_234; r11<=Pix_235; r12<=Pix_236; r13<=Pix_237; r14<=Pix_238; r15<=Pix_239; r16<=Pix_240; r17<=Pix_241; r18<=Pix_242; r19<=Pix_243; r20<=Pix_244; r21<=Pix_245; r22<=Pix_246; r23<=Pix_247; r24<=Pix_248; r25<=Pix_249; r26<=Pix_250; r27<=Pix_251; r28<=Pix_252; r29<=Pix_253; r30<=Pix_254; r31<=Pix_255; r32<=Pix_256; r33<=Pix_257; r34<=Pix_258; r35<=Pix_259; r36<=Pix_260; r37<=Pix_261; r38<=Pix_262; r39<=Pix_263; r40<=Pix_264; r41<=Pix_265; r42<=Pix_266; r43<=Pix_267; r44<=Pix_268; r45<=Pix_269; r46<=Pix_270; r47<=Pix_271; r48<=Pix_272; r49<=Pix_273; r50<=Pix_274; r51<=Pix_275; r52<=Pix_276; r53<=Pix_277; r54<=Pix_278; r55<=Pix_279; 
						select<=select+1;
					end
				8'd141:
					begin
						wr0<=w_9_280; wr1<=w_9_281; wr2<=w_9_282; wr3<=w_9_283; wr4<=w_9_284; wr5<=w_9_285; wr6<=w_9_286; wr7<=w_9_287; wr8<=w_9_288; wr9<=w_9_289; wr10<=w_9_290; wr11<=w_9_291; wr12<=w_9_292; wr13<=w_9_293; wr14<=w_9_294; wr15<=w_9_295; wr16<=w_9_296; wr17<=w_9_297; wr18<=w_9_298; wr19<=w_9_299; wr20<=w_9_300; wr21<=w_9_301; wr22<=w_9_302; wr23<=w_9_303; wr24<=w_9_304; wr25<=w_9_305; wr26<=w_9_306; wr27<=w_9_307; wr28<=w_9_308; wr29<=w_9_309; wr30<=w_9_310; wr31<=w_9_311; wr32<=w_9_312; wr33<=w_9_313; wr34<=w_9_314; wr35<=w_9_315; wr36<=w_9_316; wr37<=w_9_317; wr38<=w_9_318; wr39<=w_9_319; wr40<=w_9_320; wr41<=w_9_321; wr42<=w_9_322; wr43<=w_9_323; wr44<=w_9_324; wr45<=w_9_325; wr46<=w_9_326; wr47<=w_9_327; wr48<=w_9_328; wr49<=w_9_329; wr50<=w_9_330; wr51<=w_9_331; wr52<=w_9_332; wr53<=w_9_333; wr54<=w_9_334; wr55<=w_9_335; 
						r0<=Pix_280; r1<=Pix_281; r2<=Pix_282; r3<=Pix_283; r4<=Pix_284; r5<=Pix_285; r6<=Pix_286; r7<=Pix_287; r8<=Pix_288; r9<=Pix_289; r10<=Pix_290; r11<=Pix_291; r12<=Pix_292; r13<=Pix_293; r14<=Pix_294; r15<=Pix_295; r16<=Pix_296; r17<=Pix_297; r18<=Pix_298; r19<=Pix_299; r20<=Pix_300; r21<=Pix_301; r22<=Pix_302; r23<=Pix_303; r24<=Pix_304; r25<=Pix_305; r26<=Pix_306; r27<=Pix_307; r28<=Pix_308; r29<=Pix_309; r30<=Pix_310; r31<=Pix_311; r32<=Pix_312; r33<=Pix_313; r34<=Pix_314; r35<=Pix_315; r36<=Pix_316; r37<=Pix_317; r38<=Pix_318; r39<=Pix_319; r40<=Pix_320; r41<=Pix_321; r42<=Pix_322; r43<=Pix_323; r44<=Pix_324; r45<=Pix_325; r46<=Pix_326; r47<=Pix_327; r48<=Pix_328; r49<=Pix_329; r50<=Pix_330; r51<=Pix_331; r52<=Pix_332; r53<=Pix_333; r54<=Pix_334; r55<=Pix_335; 
						select<=select+1;
					end
				8'd142:
					begin
						wr0<=w_9_336; wr1<=w_9_337; wr2<=w_9_338; wr3<=w_9_339; wr4<=w_9_340; wr5<=w_9_341; wr6<=w_9_342; wr7<=w_9_343; wr8<=w_9_344; wr9<=w_9_345; wr10<=w_9_346; wr11<=w_9_347; wr12<=w_9_348; wr13<=w_9_349; wr14<=w_9_350; wr15<=w_9_351; wr16<=w_9_352; wr17<=w_9_353; wr18<=w_9_354; wr19<=w_9_355; wr20<=w_9_356; wr21<=w_9_357; wr22<=w_9_358; wr23<=w_9_359; wr24<=w_9_360; wr25<=w_9_361; wr26<=w_9_362; wr27<=w_9_363; wr28<=w_9_364; wr29<=w_9_365; wr30<=w_9_366; wr31<=w_9_367; wr32<=w_9_368; wr33<=w_9_369; wr34<=w_9_370; wr35<=w_9_371; wr36<=w_9_372; wr37<=w_9_373; wr38<=w_9_374; wr39<=w_9_375; wr40<=w_9_376; wr41<=w_9_377; wr42<=w_9_378; wr43<=w_9_379; wr44<=w_9_380; wr45<=w_9_381; wr46<=w_9_382; wr47<=w_9_383; wr48<=w_9_384; wr49<=w_9_385; wr50<=w_9_386; wr51<=w_9_387; wr52<=w_9_388; wr53<=w_9_389; wr54<=w_9_390; wr55<=w_9_391; 
						r0<=Pix_336; r1<=Pix_337; r2<=Pix_338; r3<=Pix_339; r4<=Pix_340; r5<=Pix_341; r6<=Pix_342; r7<=Pix_343; r8<=Pix_344; r9<=Pix_345; r10<=Pix_346; r11<=Pix_347; r12<=Pix_348; r13<=Pix_349; r14<=Pix_350; r15<=Pix_351; r16<=Pix_352; r17<=Pix_353; r18<=Pix_354; r19<=Pix_355; r20<=Pix_356; r21<=Pix_357; r22<=Pix_358; r23<=Pix_359; r24<=Pix_360; r25<=Pix_361; r26<=Pix_362; r27<=Pix_363; r28<=Pix_364; r29<=Pix_365; r30<=Pix_366; r31<=Pix_367; r32<=Pix_368; r33<=Pix_369; r34<=Pix_370; r35<=Pix_371; r36<=Pix_372; r37<=Pix_373; r38<=Pix_374; r39<=Pix_375; r40<=Pix_376; r41<=Pix_377; r42<=Pix_378; r43<=Pix_379; r44<=Pix_380; r45<=Pix_381; r46<=Pix_382; r47<=Pix_383; r48<=Pix_384; r49<=Pix_385; r50<=Pix_386; r51<=Pix_387; r52<=Pix_388; r53<=Pix_389; r54<=Pix_390; r55<=Pix_391; 
						select<=select+1;
					end
				8'd143:
					begin
						wr0<=w_9_392; wr1<=w_9_393; wr2<=w_9_394; wr3<=w_9_395; wr4<=w_9_396; wr5<=w_9_397; wr6<=w_9_398; wr7<=w_9_399; wr8<=w_9_400; wr9<=w_9_401; wr10<=w_9_402; wr11<=w_9_403; wr12<=w_9_404; wr13<=w_9_405; wr14<=w_9_406; wr15<=w_9_407; wr16<=w_9_408; wr17<=w_9_409; wr18<=w_9_410; wr19<=w_9_411; wr20<=w_9_412; wr21<=w_9_413; wr22<=w_9_414; wr23<=w_9_415; wr24<=w_9_416; wr25<=w_9_417; wr26<=w_9_418; wr27<=w_9_419; wr28<=w_9_420; wr29<=w_9_421; wr30<=w_9_422; wr31<=w_9_423; wr32<=w_9_424; wr33<=w_9_425; wr34<=w_9_426; wr35<=w_9_427; wr36<=w_9_428; wr37<=w_9_429; wr38<=w_9_430; wr39<=w_9_431; wr40<=w_9_432; wr41<=w_9_433; wr42<=w_9_434; wr43<=w_9_435; wr44<=w_9_436; wr45<=w_9_437; wr46<=w_9_438; wr47<=w_9_439; wr48<=w_9_440; wr49<=w_9_441; wr50<=w_9_442; wr51<=w_9_443; wr52<=w_9_444; wr53<=w_9_445; wr54<=w_9_446; wr55<=w_9_447; 
						r0<=Pix_392; r1<=Pix_393; r2<=Pix_394; r3<=Pix_395; r4<=Pix_396; r5<=Pix_397; r6<=Pix_398; r7<=Pix_399; r8<=Pix_400; r9<=Pix_401; r10<=Pix_402; r11<=Pix_403; r12<=Pix_404; r13<=Pix_405; r14<=Pix_406; r15<=Pix_407; r16<=Pix_408; r17<=Pix_409; r18<=Pix_410; r19<=Pix_411; r20<=Pix_412; r21<=Pix_413; r22<=Pix_414; r23<=Pix_415; r24<=Pix_416; r25<=Pix_417; r26<=Pix_418; r27<=Pix_419; r28<=Pix_420; r29<=Pix_421; r30<=Pix_422; r31<=Pix_423; r32<=Pix_424; r33<=Pix_425; r34<=Pix_426; r35<=Pix_427; r36<=Pix_428; r37<=Pix_429; r38<=Pix_430; r39<=Pix_431; r40<=Pix_432; r41<=Pix_433; r42<=Pix_434; r43<=Pix_435; r44<=Pix_436; r45<=Pix_437; r46<=Pix_438; r47<=Pix_439; r48<=Pix_440; r49<=Pix_441; r50<=Pix_442; r51<=Pix_443; r52<=Pix_444; r53<=Pix_445; r54<=Pix_446; r55<=Pix_447; 
						select<=select+1;
					end
				8'd144:
					begin
						wr0<=w_9_448; wr1<=w_9_449; wr2<=w_9_450; wr3<=w_9_451; wr4<=w_9_452; wr5<=w_9_453; wr6<=w_9_454; wr7<=w_9_455; wr8<=w_9_456; wr9<=w_9_457; wr10<=w_9_458; wr11<=w_9_459; wr12<=w_9_460; wr13<=w_9_461; wr14<=w_9_462; wr15<=w_9_463; wr16<=w_9_464; wr17<=w_9_465; wr18<=w_9_466; wr19<=w_9_467; wr20<=w_9_468; wr21<=w_9_469; wr22<=w_9_470; wr23<=w_9_471; wr24<=w_9_472; wr25<=w_9_473; wr26<=w_9_474; wr27<=w_9_475; wr28<=w_9_476; wr29<=w_9_477; wr30<=w_9_478; wr31<=w_9_479; wr32<=w_9_480; wr33<=w_9_481; wr34<=w_9_482; wr35<=w_9_483; wr36<=w_9_484; wr37<=w_9_485; wr38<=w_9_486; wr39<=w_9_487; wr40<=w_9_488; wr41<=w_9_489; wr42<=w_9_490; wr43<=w_9_491; wr44<=w_9_492; wr45<=w_9_493; wr46<=w_9_494; wr47<=w_9_495; wr48<=w_9_496; wr49<=w_9_497; wr50<=w_9_498; wr51<=w_9_499; wr52<=w_9_500; wr53<=w_9_501; wr54<=w_9_502; wr55<=w_9_503; 
						r0<=Pix_448; r1<=Pix_449; r2<=Pix_450; r3<=Pix_451; r4<=Pix_452; r5<=Pix_453; r6<=Pix_454; r7<=Pix_455; r8<=Pix_456; r9<=Pix_457; r10<=Pix_458; r11<=Pix_459; r12<=Pix_460; r13<=Pix_461; r14<=Pix_462; r15<=Pix_463; r16<=Pix_464; r17<=Pix_465; r18<=Pix_466; r19<=Pix_467; r20<=Pix_468; r21<=Pix_469; r22<=Pix_470; r23<=Pix_471; r24<=Pix_472; r25<=Pix_473; r26<=Pix_474; r27<=Pix_475; r28<=Pix_476; r29<=Pix_477; r30<=Pix_478; r31<=Pix_479; r32<=Pix_480; r33<=Pix_481; r34<=Pix_482; r35<=Pix_483; r36<=Pix_484; r37<=Pix_485; r38<=Pix_486; r39<=Pix_487; r40<=Pix_488; r41<=Pix_489; r42<=Pix_490; r43<=Pix_491; r44<=Pix_492; r45<=Pix_493; r46<=Pix_494; r47<=Pix_495; r48<=Pix_496; r49<=Pix_497; r50<=Pix_498; r51<=Pix_499; r52<=Pix_500; r53<=Pix_501; r54<=Pix_502; r55<=Pix_503; 
						select<=select+1;
					end
				8'd145:
					begin
						wr0<=w_9_504; wr1<=w_9_505; wr2<=w_9_506; wr3<=w_9_507; wr4<=w_9_508; wr5<=w_9_509; wr6<=w_9_510; wr7<=w_9_511; wr8<=w_9_512; wr9<=w_9_513; wr10<=w_9_514; wr11<=w_9_515; wr12<=w_9_516; wr13<=w_9_517; wr14<=w_9_518; wr15<=w_9_519; wr16<=w_9_520; wr17<=w_9_521; wr18<=w_9_522; wr19<=w_9_523; wr20<=w_9_524; wr21<=w_9_525; wr22<=w_9_526; wr23<=w_9_527; wr24<=w_9_528; wr25<=w_9_529; wr26<=w_9_530; wr27<=w_9_531; wr28<=w_9_532; wr29<=w_9_533; wr30<=w_9_534; wr31<=w_9_535; wr32<=w_9_536; wr33<=w_9_537; wr34<=w_9_538; wr35<=w_9_539; wr36<=w_9_540; wr37<=w_9_541; wr38<=w_9_542; wr39<=w_9_543; wr40<=w_9_544; wr41<=w_9_545; wr42<=w_9_546; wr43<=w_9_547; wr44<=w_9_548; wr45<=w_9_549; wr46<=w_9_550; wr47<=w_9_551; wr48<=w_9_552; wr49<=w_9_553; wr50<=w_9_554; wr51<=w_9_555; wr52<=w_9_556; wr53<=w_9_557; wr54<=w_9_558; wr55<=w_9_559; 
						r0<=Pix_504; r1<=Pix_505; r2<=Pix_506; r3<=Pix_507; r4<=Pix_508; r5<=Pix_509; r6<=Pix_510; r7<=Pix_511; r8<=Pix_512; r9<=Pix_513; r10<=Pix_514; r11<=Pix_515; r12<=Pix_516; r13<=Pix_517; r14<=Pix_518; r15<=Pix_519; r16<=Pix_520; r17<=Pix_521; r18<=Pix_522; r19<=Pix_523; r20<=Pix_524; r21<=Pix_525; r22<=Pix_526; r23<=Pix_527; r24<=Pix_528; r25<=Pix_529; r26<=Pix_530; r27<=Pix_531; r28<=Pix_532; r29<=Pix_533; r30<=Pix_534; r31<=Pix_535; r32<=Pix_536; r33<=Pix_537; r34<=Pix_538; r35<=Pix_539; r36<=Pix_540; r37<=Pix_541; r38<=Pix_542; r39<=Pix_543; r40<=Pix_544; r41<=Pix_545; r42<=Pix_546; r43<=Pix_547; r44<=Pix_548; r45<=Pix_549; r46<=Pix_550; r47<=Pix_551; r48<=Pix_552; r49<=Pix_553; r50<=Pix_554; r51<=Pix_555; r52<=Pix_556; r53<=Pix_557; r54<=Pix_558; r55<=Pix_559; 
						select<=select+1;
					end
				8'd146:
					begin
						wr0<=w_9_560; wr1<=w_9_561; wr2<=w_9_562; wr3<=w_9_563; wr4<=w_9_564; wr5<=w_9_565; wr6<=w_9_566; wr7<=w_9_567; wr8<=w_9_568; wr9<=w_9_569; wr10<=w_9_570; wr11<=w_9_571; wr12<=w_9_572; wr13<=w_9_573; wr14<=w_9_574; wr15<=w_9_575; wr16<=w_9_576; wr17<=w_9_577; wr18<=w_9_578; wr19<=w_9_579; wr20<=w_9_580; wr21<=w_9_581; wr22<=w_9_582; wr23<=w_9_583; wr24<=w_9_584; wr25<=w_9_585; wr26<=w_9_586; wr27<=w_9_587; wr28<=w_9_588; wr29<=w_9_589; wr30<=w_9_590; wr31<=w_9_591; wr32<=w_9_592; wr33<=w_9_593; wr34<=w_9_594; wr35<=w_9_595; wr36<=w_9_596; wr37<=w_9_597; wr38<=w_9_598; wr39<=w_9_599; wr40<=w_9_600; wr41<=w_9_601; wr42<=w_9_602; wr43<=w_9_603; wr44<=w_9_604; wr45<=w_9_605; wr46<=w_9_606; wr47<=w_9_607; wr48<=w_9_608; wr49<=w_9_609; wr50<=w_9_610; wr51<=w_9_611; wr52<=w_9_612; wr53<=w_9_613; wr54<=w_9_614; wr55<=w_9_615; 
						r0<=Pix_560; r1<=Pix_561; r2<=Pix_562; r3<=Pix_563; r4<=Pix_564; r5<=Pix_565; r6<=Pix_566; r7<=Pix_567; r8<=Pix_568; r9<=Pix_569; r10<=Pix_570; r11<=Pix_571; r12<=Pix_572; r13<=Pix_573; r14<=Pix_574; r15<=Pix_575; r16<=Pix_576; r17<=Pix_577; r18<=Pix_578; r19<=Pix_579; r20<=Pix_580; r21<=Pix_581; r22<=Pix_582; r23<=Pix_583; r24<=Pix_584; r25<=Pix_585; r26<=Pix_586; r27<=Pix_587; r28<=Pix_588; r29<=Pix_589; r30<=Pix_590; r31<=Pix_591; r32<=Pix_592; r33<=Pix_593; r34<=Pix_594; r35<=Pix_595; r36<=Pix_596; r37<=Pix_597; r38<=Pix_598; r39<=Pix_599; r40<=Pix_600; r41<=Pix_601; r42<=Pix_602; r43<=Pix_603; r44<=Pix_604; r45<=Pix_605; r46<=Pix_606; r47<=Pix_607; r48<=Pix_608; r49<=Pix_609; r50<=Pix_610; r51<=Pix_611; r52<=Pix_612; r53<=Pix_613; r54<=Pix_614; r55<=Pix_615; 
						select<=select+1;
					end
				8'd147:
					begin
						wr0<=w_9_616; wr1<=w_9_617; wr2<=w_9_618; wr3<=w_9_619; wr4<=w_9_620; wr5<=w_9_621; wr6<=w_9_622; wr7<=w_9_623; wr8<=w_9_624; wr9<=w_9_625; wr10<=w_9_626; wr11<=w_9_627; wr12<=w_9_628; wr13<=w_9_629; wr14<=w_9_630; wr15<=w_9_631; wr16<=w_9_632; wr17<=w_9_633; wr18<=w_9_634; wr19<=w_9_635; wr20<=w_9_636; wr21<=w_9_637; wr22<=w_9_638; wr23<=w_9_639; wr24<=w_9_640; wr25<=w_9_641; wr26<=w_9_642; wr27<=w_9_643; wr28<=w_9_644; wr29<=w_9_645; wr30<=w_9_646; wr31<=w_9_647; wr32<=w_9_648; wr33<=w_9_649; wr34<=w_9_650; wr35<=w_9_651; wr36<=w_9_652; wr37<=w_9_653; wr38<=w_9_654; wr39<=w_9_655; wr40<=w_9_656; wr41<=w_9_657; wr42<=w_9_658; wr43<=w_9_659; wr44<=w_9_660; wr45<=w_9_661; wr46<=w_9_662; wr47<=w_9_663; wr48<=w_9_664; wr49<=w_9_665; wr50<=w_9_666; wr51<=w_9_667; wr52<=w_9_668; wr53<=w_9_669; wr54<=w_9_670; wr55<=w_9_671; 
						r0<=Pix_616; r1<=Pix_617; r2<=Pix_618; r3<=Pix_619; r4<=Pix_620; r5<=Pix_621; r6<=Pix_622; r7<=Pix_623; r8<=Pix_624; r9<=Pix_625; r10<=Pix_626; r11<=Pix_627; r12<=Pix_628; r13<=Pix_629; r14<=Pix_630; r15<=Pix_631; r16<=Pix_632; r17<=Pix_633; r18<=Pix_634; r19<=Pix_635; r20<=Pix_636; r21<=Pix_637; r22<=Pix_638; r23<=Pix_639; r24<=Pix_640; r25<=Pix_641; r26<=Pix_642; r27<=Pix_643; r28<=Pix_644; r29<=Pix_645; r30<=Pix_646; r31<=Pix_647; r32<=Pix_648; r33<=Pix_649; r34<=Pix_650; r35<=Pix_651; r36<=Pix_652; r37<=Pix_653; r38<=Pix_654; r39<=Pix_655; r40<=Pix_656; r41<=Pix_657; r42<=Pix_658; r43<=Pix_659; r44<=Pix_660; r45<=Pix_661; r46<=Pix_662; r47<=Pix_663; r48<=Pix_664; r49<=Pix_665; r50<=Pix_666; r51<=Pix_667; r52<=Pix_668; r53<=Pix_669; r54<=Pix_670; r55<=Pix_671; 
						select<=select+1;
					end
				8'd148:
					begin
						wr0<=w_9_672; wr1<=w_9_673; wr2<=w_9_674; wr3<=w_9_675; wr4<=w_9_676; wr5<=w_9_677; wr6<=w_9_678; wr7<=w_9_679; wr8<=w_9_680; wr9<=w_9_681; wr10<=w_9_682; wr11<=w_9_683; wr12<=w_9_684; wr13<=w_9_685; wr14<=w_9_686; wr15<=w_9_687; wr16<=w_9_688; wr17<=w_9_689; wr18<=w_9_690; wr19<=w_9_691; wr20<=w_9_692; wr21<=w_9_693; wr22<=w_9_694; wr23<=w_9_695; wr24<=w_9_696; wr25<=w_9_697; wr26<=w_9_698; wr27<=w_9_699; wr28<=w_9_700; wr29<=w_9_701; wr30<=w_9_702; wr31<=w_9_703; wr32<=w_9_704; wr33<=w_9_705; wr34<=w_9_706; wr35<=w_9_707; wr36<=w_9_708; wr37<=w_9_709; wr38<=w_9_710; wr39<=w_9_711; wr40<=w_9_712; wr41<=w_9_713; wr42<=w_9_714; wr43<=w_9_715; wr44<=w_9_716; wr45<=w_9_717; wr46<=w_9_718; wr47<=w_9_719; wr48<=w_9_720; wr49<=w_9_721; wr50<=w_9_722; wr51<=w_9_723; wr52<=w_9_724; wr53<=w_9_725; wr54<=w_9_726; wr55<=w_9_727; 
						r0<=Pix_672; r1<=Pix_673; r2<=Pix_674; r3<=Pix_675; r4<=Pix_676; r5<=Pix_677; r6<=Pix_678; r7<=Pix_679; r8<=Pix_680; r9<=Pix_681; r10<=Pix_682; r11<=Pix_683; r12<=Pix_684; r13<=Pix_685; r14<=Pix_686; r15<=Pix_687; r16<=Pix_688; r17<=Pix_689; r18<=Pix_690; r19<=Pix_691; r20<=Pix_692; r21<=Pix_693; r22<=Pix_694; r23<=Pix_695; r24<=Pix_696; r25<=Pix_697; r26<=Pix_698; r27<=Pix_699; r28<=Pix_700; r29<=Pix_701; r30<=Pix_702; r31<=Pix_703; r32<=Pix_704; r33<=Pix_705; r34<=Pix_706; r35<=Pix_707; r36<=Pix_708; r37<=Pix_709; r38<=Pix_710; r39<=Pix_711; r40<=Pix_712; r41<=Pix_713; r42<=Pix_714; r43<=Pix_715; r44<=Pix_716; r45<=Pix_717; r46<=Pix_718; r47<=Pix_719; r48<=Pix_720; r49<=Pix_721; r50<=Pix_722; r51<=Pix_723; r52<=Pix_724; r53<=Pix_725; r54<=Pix_726; r55<=Pix_727; 
						select<=select+1;
					end
				8'd149:
					begin
						wr0<=w_9_728; wr1<=w_9_729; wr2<=w_9_730; wr3<=w_9_731; wr4<=w_9_732; wr5<=w_9_733; wr6<=w_9_734; wr7<=w_9_735; wr8<=w_9_736; wr9<=w_9_737; wr10<=w_9_738; wr11<=w_9_739; wr12<=w_9_740; wr13<=w_9_741; wr14<=w_9_742; wr15<=w_9_743; wr16<=w_9_744; wr17<=w_9_745; wr18<=w_9_746; wr19<=w_9_747; wr20<=w_9_748; wr21<=w_9_749; wr22<=w_9_750; wr23<=w_9_751; wr24<=w_9_752; wr25<=w_9_753; wr26<=w_9_754; wr27<=w_9_755; wr28<=w_9_756; wr29<=w_9_757; wr30<=w_9_758; wr31<=w_9_759; wr32<=w_9_760; wr33<=w_9_761; wr34<=w_9_762; wr35<=w_9_763; wr36<=w_9_764; wr37<=w_9_765; wr38<=w_9_766; wr39<=w_9_767; wr40<=w_9_768; wr41<=w_9_769; wr42<=w_9_770; wr43<=w_9_771; wr44<=w_9_772; wr45<=w_9_773; wr46<=w_9_774; wr47<=w_9_775; wr48<=w_9_776; wr49<=w_9_777; wr50<=w_9_778; wr51<=w_9_779; wr52<=w_9_780; wr53<=w_9_781; wr54<=w_9_782; wr55<=w_9_783; 
						r0<=Pix_728; r1<=Pix_729; r2<=Pix_730; r3<=Pix_731; r4<=Pix_732; r5<=Pix_733; r6<=Pix_734; r7<=Pix_735; r8<=Pix_736; r9<=Pix_737; r10<=Pix_738; r11<=Pix_739; r12<=Pix_740; r13<=Pix_741; r14<=Pix_742; r15<=Pix_743; r16<=Pix_744; r17<=Pix_745; r18<=Pix_746; r19<=Pix_747; r20<=Pix_748; r21<=Pix_749; r22<=Pix_750; r23<=Pix_751; r24<=Pix_752; r25<=Pix_753; r26<=Pix_754; r27<=Pix_755; r28<=Pix_756; r29<=Pix_757; r30<=Pix_758; r31<=Pix_759; r32<=Pix_760; r33<=Pix_761; r34<=Pix_762; r35<=Pix_763; r36<=Pix_764; r37<=Pix_765; r38<=Pix_766; r39<=Pix_767; r40<=Pix_768; r41<=Pix_769; r42<=Pix_770; r43<=Pix_771; r44<=Pix_772; r45<=Pix_773; r46<=Pix_774; r47<=Pix_775; r48<=Pix_776; r49<=Pix_777; r50<=Pix_778; r51<=Pix_779; r52<=Pix_780; r53<=Pix_781; r54<=Pix_782; r55<=Pix_783; 
						select<=select+1;
					end
				8'd150:
					begin
						bias_p<=px_784;
						bias_w<=w_9_784;
						select<=8'd0;
					end

				//************** finish off
				//need 8 more extra cycle;
			default: select<=8'bxxxxxxxx; 
			endcase	
		end
	end	
	
always @(posedge clk or negedge GlobalReset) begin
	if ((GlobalReset == 1'b0))
		begin
			//counter <= {(6){1'b0}};
			state<={(6){1'b0}};
			//neuron_flag<={(4){1'b0}};
			flag_1st<=0;
		
			//seq <= {(8){1'b0}};
			//reset all the register //not done
		end
	else
		begin
			case(state)
			
				6'd0: 
				begin
					state<=state+1;
				end
				6'd1: 
				begin
					state<=state+1;
				end
				6'd2: 
				begin
					state<=state+1;
				end
				6'd3: 
				begin
					state<=state+1;
				end
				6'd4: 
				begin
					state<=state+1;
				end
				6'd5: 
				begin
					state<=state+1;
				end
				6'd6: 
				begin
					state<=state+1;
				end
				6'd7: 
				begin
					state<=state+1;
				end
				6'd8: 
				begin
					state<=state+1;
				end
				6'd9: 
				begin
					state<=state+1;
				end
				6'd10: 
				begin
					state<=state+1;
				end
				6'd11: 
				begin
					state<=state+1;
				end
				6'd12: 
				begin
					state<=state+1;
				end
				6'd13: 
				begin
					state<=state+1;
				end
				6'd14: 
				begin
					state<=state+1;
				end
				6'd15: 
				begin
					state<=state+1;
				end
				6'd16: 
				begin
					state<=state+1;
				end
				6'd17: 
				begin
					state<=state+1;
				end
				6'd18: 
				begin
					state<=state+1;
				end
				6'd19: 
				begin
					state<=6'd35;
				end				
					/*counter<=counter+1;
					if (counter==6'd20) 
					begin
						//out_0<=out_7th_temp;
						state<=8'd15;
						counter<=0;
						//$display(out_0);
					end
					else
					begin
						state<=6'd0;
					end*/
					
				6'd20:
				begin				
					//counter<=counter+1;
					out_1<=out_7th_temp;
					state<=state+1; 
					//$display(out_1);					
				end
				6'd21:
				begin
					//counter<=counter+1;
					out_2<=out_7th_temp;
					state<=state+1;
					
				end
				6'd22:
				begin
					//counter<=counter+1;
					out_3<=out_7th_temp;
					state<=state+1;

				end
				6'd23: 
				begin	
					//counter<=counter+1;
					out_4<=out_7th_temp;
					state<=state+1; 			
				end
				6'd24: 
				begin	
					//counter<=counter+1;
					out_5<=out_7th_temp;
					state<=state+1;
					//$display("5");
					//$display(out_5);					
				end
				6'd25:
				begin
					//counter<=counter+1;
					out_6<=out_7th_temp;
					state<=state+1; 
				end
				6'd26: 
				begin	
					//counter<=counter+1;
					out_7<=out_7th_temp;
					state<=state+1; 
				end
				6'd27: 
				begin	
					//counter<=counter+1;
					out_8<=out_7th_temp;
					state<=state+1; 
				end
				6'd28: 
				begin	
					//counter<=counter+1;
					out_9<=out_7th_temp;
					state<=state+1; 
				end
				6'd29: 
				begin	
					//counter<=counter+1;
					out_10<=out_7th_temp;
					state<=state+1; 
				end
				6'd30: 
				begin	
					//counter<=counter+1;
					out_11<=out_7th_temp;
					state<=state+1; 
				end
				6'd31: 
				begin	
					//counter<=counter+1;
					out_12<=out_7th_temp;
					state<=state+1; 				
				end
				6'd32: 
				begin	
					//$display("enter 13th");
					//counter<=0;
					out_13<=out_7th_temp;	
					state<=state+1;//next cycle out_0 again
					flag_1st<=1;
				end	
				6'd33:
				begin
					state<=state+1;
					flag_1st<=0;//extra cycle for bias
				end
				6'd34:
				begin
					if(!flag_s)
					begin
						out_0<=out_7th_temp;
						//counter<=counter+1;
						state<=6'd20;
					end
					else
					begin
					
						state<=6'd38;
					end
				end
				6'd35: 
				begin
					state<=6'd34;
				end				

				
				6'd38:
				begin
					if(Input_Valid)
					begin
						//counter<=0;
						state<=6'd0;
					end
					else
					begin
						state<=6'd38;
					end
				
					//$display("done!");
				end
					//$display(out_0);*/
				//end
							
			default: state<=5'bxxxxx;
			endcase	
		end 

	end
always @(posedge clk or negedge GlobalReset) begin
	if (GlobalReset == 1'b0)
		begin
		//reset
		status<=0;
		//sum_cnt<=0;
		flagging_neuron<=0;
		flag_stop<=0;
		ov<=0;
		end
	else
		begin
			case(status)
				5'd0:
				begin
				      ov<=0;
					  flagging_neuron<=0;
					  if(flag_1st)
					  begin
						//sum_cnt<=0;
						status<=status+1;
					  end
					  else
					  begin
						status<=5'd0;
						//ov<=0;
					  end
				end	  
				
				5'd1:
				begin
					status<=status+1;
				end
				5'd2:
				begin
					status<=status+1;
				end
				5'd3:
				begin
					status<=status+1;
				end
				5'd4:
				begin
					status<=status+1;
				end
				5'd5:
				begin
					status<=status+1;
				end
				5'd6:
				begin
					status<=status+1;
				end
				5'd7:
				begin
					status<=status+1;
				end
				5'd8:
				begin
					status<=status+2;
				end
				
				5'd10:
				begin
					/*if (sum_cnt>8)
					begin*/
					if(!flag_s)
					begin
					flagging_neuron<=1;
					status<=5'd0;
					flag_stop<=1;
					end
					else
					begin
					
					status<=5'd11;
					end
						
						
	
				
				end
				
				5'd11:
					begin
						if(!flag_stop)
						begin	
						status<=5'd0;
						
						end
						else
						begin
							buffer0<=out_total_0;
							buffer1<=out_total_1;
							buffer2<=out_total_2;   
							buffer3<=out_total_3;
							buffer4<=out_total_4;
							buffer5<=out_total_5;
							buffer6<=out_total_6;
							buffer7<=out_total_7;
							buffer8<=out_total_8;
							buffer9<=out_total_9;
							status<=status+1;
	
						end
					end
				
				5'd12:
					begin
						if(buffer0[25])
						begin	
							buffer0<=0;
						end
						if (buffer1[25])
						begin		
							buffer1<=0;
						end
						if (buffer2[25])
						begin		
							buffer2<=0;
						end	
						if (buffer3[25])
						begin		
							buffer3<=0;
						end	
						if (buffer4[25])
						begin		
							buffer4<=0;
						end	
						if (buffer5[25])
						begin		
							buffer5<=0;
						end	
						if (buffer6[25])
						begin		
							buffer6<=0;
						end	
						if (buffer7[25])
						begin		
							buffer7<=0;
						end	
						if (buffer8[25])
						begin		
							buffer8<=0;
						end
						if (buffer9[25])
						begin		
							buffer9<=0;
						end							
						else
						begin
							
						end
						status<=status+1;
						/*if (buffer0 < buffer1)
						begin	
							buffer5 <= buffer1;
						end
						else
						begin
							buffer5 <= buffer0;
						end
						if (buffer2 < buffer3)
						begin	
							buffer6 <= buffer3;
						end
						else
						begin
							buffer6 <= buffer2;
						end	
						status<=8'd4;*/
					end
				5'd13:
					begin	
						if(buffer0<buffer1)
						begin
						temp_buffer0<=buffer1;
						end
						else
						begin
						temp_buffer0<=buffer0;
						end
						if(buffer2<buffer3)
						begin
						temp_buffer1<=buffer3;
						end
						else
						begin
						temp_buffer1<=buffer2;
						end
						if(buffer4<buffer5)
						begin
						temp_buffer2<=buffer5;
						end
						else
						begin
						temp_buffer2<=buffer4;
						end
						if(buffer6<buffer7)
						begin
						temp_buffer3<=buffer7;
						end
						else
						begin
						temp_buffer3<=buffer6;
						end
						if(buffer8<buffer9)
						begin
						temp_buffer4<=buffer9;
						end
						else
						begin
						temp_buffer4<=buffer8;
						end						
						status<=status+1;
					end
				
				5'd14:		
					begin
						if (temp_buffer0< temp_buffer1)
						begin		
							temp_buffer5 <= temp_buffer1;
						end
						else
						begin
							temp_buffer5 <= temp_buffer0;
						end
						if (temp_buffer2< temp_buffer3)
						begin		
							temp_buffer6 <= temp_buffer3;
						end
						else
						begin
							temp_buffer6 <= temp_buffer2;
						end
						
				
						status<=status+1;
					end		// Get the answer
				5'd15:
					begin
						if (temp_buffer4< temp_buffer5)
						begin		
							temp_buffer7 <= temp_buffer5;
						end
						else
						begin
							temp_buffer7 <= temp_buffer4;
						end
						status<=status+1;
					
					end
				5'd16:
					begin
						if (temp_buffer6< temp_buffer7)
						begin		
							buffer_select <= temp_buffer7;
						end
						else
						begin
							buffer_select <= temp_buffer6;
						end
						buff<=1;
						status<=status+1;
					end
				
				5'd17:
					begin	
						
						
						ov<=1;
						buff<=0;
						
						flag_stop<=0;
						//flag_1st<=0;
						//neuron_flag<=0;
						//sum_cnt<=0;
						status<=5'd0;
			

					
					end

					
					
				default:status<=4'bxxxx;
					
			
			
			
			
			
			endcase
		end

end
always @(posedge clk or negedge GlobalReset) begin
	if ((GlobalReset == 1'b0))
		begin
			flag_s<=0;
			//flagging_neuron<=0;
			neuron_flag<=0;
		end	
	else
	begin
		if(Input_Valid)
		begin
			flag_s<=0;
		end
		else
		begin
		end
			case(neuron_flag)
				4'd0:
				begin
					if(flagging_neuron)
					begin
						out_total_0<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else					
						neuron_flag<=4'd0;					//$display("This is out total 0");
				end
				4'd1:
				begin

					if(flagging_neuron)
					begin
						out_total_1<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else
					begin
						neuron_flag<=4'd1;	
					end					
										//$display("This is out total 1");
				end
				4'd2:
				begin
										
					if(flagging_neuron)
					begin
						out_total_2<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else	
					begin
						neuron_flag<=4'd2;	//out_total_2<=temp_output;
					end					//$display("This is out total 2");
				end
				4'd3:
				begin						
					if(flagging_neuron)
					begin
						out_total_3<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else
					begin
						neuron_flag<=4'd3;
					end					//status<=5'd0;
			
										
										//$display("This is out total 3");
				end
				4'd4:
				begin

					if(flagging_neuron)
					begin
						out_total_4<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else
					begin
						neuron_flag<=4'd4;
					end					//$display("This is out total 4");
				end
				4'd5:
				begin
					if(flagging_neuron)
					begin
						out_total_5<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else
					begin
						neuron_flag<=4'd5;
					end					//status<=5'd0;

				//$display("This is out total 5");
				end						 
				4'd6:
				begin
					if(flagging_neuron)
					begin
						out_total_6<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else	
					begin
						neuron_flag<=4'd6;
					end					//$display("This is out total 6");
				end
				4'd7:
				begin
					if(flagging_neuron)
					begin
						out_total_7<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else	
					begin
						neuron_flag<=4'd7;
					end		
				end
				4'd8:
					if(flagging_neuron)
					begin
						out_total_8<=temp_output;
						neuron_flag<=neuron_flag+1;
						//flagging_neuron<=0;
					end
					//status<=5'd0;
					else	
					begin
						neuron_flag<=4'd8;
					end	
				4'd9:
					begin
										
						if(flagging_neuron)
						begin
							out_total_9<=temp_output;
							neuron_flag<=0;
							//flagging_neuron<=0;
							flag_s<=1;
						end
						//status<=5'd0;
						else	
						begin
							neuron_flag<=4'd9;
						end			
									
									
					end		
			default: neuron_flag<=4'bxxxx;
			endcase		
		
		
	end
end
always @(posedge clk or negedge GlobalReset) begin
	if ((GlobalReset == 1'b0))
		begin
			
	
		end	
	else
	begin
		if(buff)
		begin
			if(buffer_select==out_total_0)
				begin	
					outBuffer<=4'd0;
				end
			else if(buffer_select==out_total_1)
				begin	
						outBuffer<=4'd1;
				end
			else if(buffer_select==out_total_2)
				begin	
					outBuffer<=4'd2;
				end
			else if(buffer_select==out_total_3)
				begin	
					outBuffer<=4'd3;
				end
			else if(buffer_select==out_total_4)
				begin	
					outBuffer<=4'd4;
				end
			else if(buffer_select==out_total_5)
				begin	
					outBuffer<=4'd5;
				end
			else if(buffer_select==out_total_6)
				begin	
							outBuffer<=4'd6;
				end
			else if(buffer_select==out_total_7)
				begin	
					outBuffer<=4'd7;
				end
			else if(buffer_select==out_total_8)
				begin	
					outBuffer<=4'd8;
				end
			else if(buffer_select==out_total_9)
				begin	
					outBuffer<=4'd9;
				end
			else
				begin
					outBuffer<=4'bxxxx;
				end						
	
		end
	end
end

endmodule
							
							
					